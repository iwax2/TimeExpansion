
module b15 ( CLOCK, RESET, HOLD, NA_n, BS16_n, READY_n, BE_n, Address, W_R_n, 
        D_C_n, M_IO_n, ADS_n, Datai, Datao );
  output [3:0] BE_n;
  output [29:0] Address;
  input [31:0] Datai;
  output [31:0] Datao;
  input CLOCK, RESET, HOLD, NA_n, BS16_n, READY_n;
  output W_R_n, D_C_n, M_IO_n, ADS_n;
  wire   N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N818, N819, N1750,
         N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759, N1760,
         N1761, N1762, N1763, N1764, N2579, N2580, N2581, N2582, N2583, N2584,
         N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594,
         N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604,
         N2605, N2606, N2607, N2608, N2609, N2787, N2788, N2789, N2790, N2791,
         N2792, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, U3_U1_Z_0,
         U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3, U3_U1_Z_4, U3_U1_Z_5, U3_U1_Z_6,
         U3_U1_Z_7, U3_U1_Z_8, U3_U1_Z_9, U3_U1_Z_10, U3_U1_Z_11, U3_U1_Z_12,
         U3_U1_Z_13, U3_U1_Z_14, U3_U1_Z_15, U3_U1_Z_16, U3_U1_Z_17,
         U3_U1_Z_18, U3_U1_Z_19, U3_U1_Z_20, U3_U1_Z_21, U3_U1_Z_22,
         U3_U1_Z_23, U3_U1_Z_24, U3_U1_Z_25, U3_U1_Z_26, U3_U1_Z_27,
         U3_U1_Z_28, U3_U1_Z_29, U3_U2_Z_0, U3_U3_Z_0, U3_U3_Z_1, U3_U3_Z_2,
         U3_U3_Z_3, U3_U3_Z_4, U3_U3_Z_5, U3_U3_Z_6, U3_U3_Z_7, U3_U3_Z_8,
         U3_U3_Z_9, U3_U3_Z_10, U3_U3_Z_11, U3_U3_Z_12, U3_U3_Z_13, U3_U3_Z_14,
         U3_U4_Z_0, U3_U5_Z_0, U3_U5_Z_1, U3_U5_Z_2, U3_U5_Z_3, U3_U5_Z_4,
         U3_U5_Z_5, U3_U5_Z_6, U3_U5_Z_7, U3_U5_Z_8, U3_U5_Z_9, U3_U5_Z_10,
         U3_U5_Z_11, U3_U5_Z_12, U3_U5_Z_13, U3_U5_Z_14, U3_U5_Z_15,
         U3_U5_Z_16, U3_U5_Z_17, U3_U5_Z_18, U3_U5_Z_19, U3_U5_Z_20,
         U3_U5_Z_21, U3_U5_Z_22, U3_U5_Z_23, U3_U5_Z_24, U3_U5_Z_25,
         U3_U5_Z_26, U3_U5_Z_27, U3_U5_Z_28, U3_U5_Z_29, U3_U5_Z_30, U3_U6_Z_0,
         U3_U6_Z_1, U3_U6_Z_2, U3_U6_Z_3, U3_U6_Z_4, U3_U6_Z_5, U3_U6_Z_6,
         U3_U6_Z_7, U3_U6_Z_8, U3_U6_Z_9, U3_U6_Z_10, U3_U6_Z_11, U3_U6_Z_12,
         U3_U6_Z_13, U3_U6_Z_14, U3_U6_Z_15, U3_U6_Z_16, U3_U6_Z_17,
         U3_U6_Z_18, U3_U6_Z_19, U3_U6_Z_20, U3_U6_Z_21, U3_U6_Z_22,
         U3_U6_Z_23, U3_U6_Z_24, U3_U6_Z_25, U3_U6_Z_26, U3_U6_Z_27,
         U3_U6_Z_28, U3_U6_Z_29, U3_U6_Z_30, U3_U7_Z_0, U3_U7_Z_1, U3_U7_Z_2,
         U3_U7_Z_3, U3_U8_Z_1, U3_U8_Z_2, U3_U8_Z_3, U3_U8_Z_4, U3_U8_Z_5,
         U3_U8_Z_6, U3_U8_Z_7, U3_U13_Z_0, U3_U13_Z_1, U3_U13_Z_2, U3_U13_Z_3,
         U3_U13_Z_4, U3_U13_Z_5, U3_U13_Z_6, U3_U13_Z_7, U3_U13_Z_8,
         U3_U13_Z_9, U3_U13_Z_10, U3_U13_Z_11, U3_U13_Z_12, U3_U13_Z_13,
         U3_U13_Z_14, U3_U13_Z_15, U3_U13_Z_16, U3_U13_Z_17, U3_U13_Z_18,
         U3_U13_Z_19, U3_U13_Z_20, U3_U13_Z_21, U3_U13_Z_22, U3_U13_Z_23,
         U3_U13_Z_24, U3_U13_Z_25, U3_U13_Z_26, U3_U13_Z_27, U3_U13_Z_28,
         U3_U13_Z_29, U3_U13_Z_30, U3_U13_Z_31, U3_U14_Z_0, U3_U14_Z_1,
         U3_U14_Z_2, U3_U14_Z_3, U3_U14_Z_4, U3_U14_Z_5, U3_U14_Z_6,
         U3_U14_Z_7, U3_U18_Z_0, U3_U18_Z_1, U3_U18_Z_2, U3_U18_Z_3,
         U3_U18_Z_4, U3_U18_Z_5, U3_U18_Z_6, U3_U18_Z_7, U3_U18_Z_8,
         U3_U18_Z_9, U3_U18_Z_10, U3_U18_Z_11, U3_U18_Z_12, U3_U18_Z_13,
         U3_U18_Z_14, U3_U18_Z_15, U3_U18_Z_16, U3_U18_Z_17, U3_U18_Z_18,
         U3_U18_Z_19, U3_U18_Z_20, U3_U18_Z_21, U3_U18_Z_22, U3_U18_Z_23,
         U3_U18_Z_24, U3_U18_Z_25, U3_U18_Z_26, U3_U18_Z_27, U3_U18_Z_28,
         U3_U18_Z_29, U3_U18_Z_30, U3_U18_Z_31, U3_U19_Z_0, U3_U19_Z_2,
         U3_U19_Z_3, U3_U19_Z_4, U3_U19_Z_5, U3_U19_Z_6, U3_U19_Z_7,
         U3_U21_Z_0, U3_U21_Z_16, U3_U21_Z_17, U3_U21_Z_18, U3_U21_Z_19,
         U3_U21_Z_20, U3_U21_Z_21, U3_U21_Z_22, U3_U21_Z_23, U3_U21_Z_24,
         U3_U21_Z_25, U3_U21_Z_26, U3_U21_Z_27, U3_U21_Z_28, U3_U21_Z_29,
         U3_U21_Z_30, U3_U22_Z_0, U3_U22_Z_1, U3_U22_Z_2, U3_U22_Z_3,
         U3_U22_Z_4, U3_U22_Z_5, U3_U22_Z_6, U3_U22_Z_7, U3_U22_Z_8,
         U3_U22_Z_9, U3_U22_Z_10, U3_U22_Z_11, U3_U22_Z_12, U3_U22_Z_13,
         U3_U22_Z_14, U3_U22_Z_15, U3_U22_Z_20, U3_U22_Z_21, U3_U22_Z_22,
         U3_U22_Z_23, U3_U22_Z_24, U3_U22_Z_25, U3_U22_Z_26, U3_U22_Z_27,
         U3_U22_Z_28, U3_U22_Z_29, U3_U22_Z_30, U3_U22_Z_31, U3_U23_Z_0, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3233, n3234, n3236, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n5296, n5298,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5397, n5409, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5429, n5430, n5488, n5489, n5490, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n22, n35, n73, n567, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n3020,
         n3232, n3235, n3237, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, r1165_n17, r1165_n16, r1165_n15,
         r1165_n14, r1165_n13, r1165_n12, r1165_n11, r1165_n10, r1165_n9,
         r1165_n8, r1165_n7, r1165_n6, r1165_n5, r1165_n4, r1165_n3, r1165_n2,
         r1165_n1, r1164_n145, r1164_n144, r1164_n143, r1164_n142, r1164_n141,
         r1164_n140, r1164_n139, r1164_n138, r1164_n137, r1164_n136,
         r1164_n135, r1164_n134, r1164_n133, r1164_n132, r1164_n131,
         r1164_n130, r1164_n129, r1164_n128, r1164_n127, r1164_n126,
         r1164_n125, r1164_n124, r1164_n123, r1164_n122, r1164_n121,
         r1164_n120, r1164_n119, r1164_n118, r1164_n117, r1164_n116,
         r1164_n115, r1164_n114, r1164_n113, r1164_n112, r1164_n111,
         r1164_n110, r1164_n109, r1164_n108, r1164_n107, r1164_n106,
         r1164_n105, r1164_n104, r1164_n103, r1164_n102, r1164_n101,
         r1164_n100, r1164_n99, r1164_n98, r1164_n97, r1164_n96, r1164_n95,
         r1164_n94, r1164_n93, r1164_n92, r1164_n91, r1164_n90, r1164_n89,
         r1164_n88, r1164_n87, r1164_n86, r1164_n85, r1164_n84, r1164_n83,
         r1164_n82, r1164_n81, r1164_n80, r1164_n79, r1164_n78, r1164_n77,
         r1164_n76, r1164_n75, r1164_n74, r1164_n73, r1164_n72, r1164_n71,
         r1164_n70, r1164_n69, r1164_n68, r1164_n67, r1164_n66, r1164_n65,
         r1164_n64, r1164_n63, r1164_n62, r1164_n61, r1164_n60, r1164_n59,
         r1164_n58, r1164_n57, r1164_n56, r1164_n55, r1164_n54, r1164_n53,
         r1164_n52, r1164_n51, r1164_n50, r1164_n49, r1164_n48, r1164_n47,
         r1164_n46, r1164_n45, r1164_n44, r1164_n43, r1164_n42, r1164_n41,
         r1164_n40, r1164_n39, r1164_n38, r1164_n37, r1164_n36, r1164_n35,
         r1164_n34, r1164_n33, r1164_n32, r1164_n31, r1164_n30, r1164_n29,
         r1164_n28, r1164_n27, r1164_n26, r1164_n25, r1164_n24, r1164_n23,
         r1164_n22, r1164_n21, r1164_n20, r1164_n19, r1164_n18, r1164_n17,
         r1164_n16, r1164_n15, r1164_n14, r1164_n13, r1164_n12, r1164_n11,
         r1164_n10, r1164_n9, r1164_n8, r1164_n7, r1164_n6, r1164_n5, r1164_n4,
         r1164_n3, r1164_n2, r1164_n1, r1166_n107, r1166_n106, r1166_n105,
         r1166_n104, r1166_n103, r1166_n102, r1166_n101, r1166_n100, r1166_n99,
         r1166_n98, r1166_n97, r1166_n96, r1166_n95, r1166_n94, r1166_n93,
         r1166_n92, r1166_n91, r1166_n90, r1166_n89, r1166_n88, r1166_n87,
         r1166_n86, r1166_n85, r1166_n84, r1166_n83, r1166_n82, r1166_n81,
         r1166_n80, r1166_n79, r1166_n78, r1166_n77, r1166_n76, r1166_n75,
         r1166_n74, r1166_n73, r1166_n72, r1166_n71, r1166_n70, r1166_n69,
         r1166_n68, r1166_n67, r1166_n66, r1166_n65, r1166_n64, r1166_n63,
         r1166_n62, r1166_n61, r1166_n60, r1166_n59, r1166_n58, r1166_n57,
         r1166_n56, r1166_n55, r1166_n54, r1166_n53, r1166_n52, r1166_n51,
         r1166_n50, r1166_n49, r1166_n48, r1166_n47, r1166_n46, r1166_n45,
         r1166_n44, r1166_n43, r1166_n42, r1166_n41, r1166_n40, r1166_n39,
         r1166_n38, r1166_n37, r1166_n36, r1166_n35, r1166_n34, r1166_n33,
         r1166_n32, r1166_n31, r1166_n30, r1166_n29, r1166_n28, r1166_n27,
         r1166_n26, r1166_n25, r1166_n24, r1166_n23, r1166_n22, r1166_n21,
         r1166_n20, r1166_n19, r1166_n18, r1166_n17, r1166_n16, r1166_n15,
         r1166_n14, r1166_n13, r1166_n12, r1166_n11, r1166_n10, r1166_n9,
         r1166_n8, r1166_n7, r1166_n6, r1166_n5, r1166_n4, r1166_n3, r1166_n2,
         r1166_n1, r253_n148, r253_n147, r253_n146, r253_n145, r253_n144,
         r253_n143, r253_n142, r253_n141, r253_n140, r253_n139, r253_n138,
         r253_n137, r253_n136, r253_n135, r253_n134, r253_n133, r253_n132,
         r253_n131, r253_n130, r253_n129, r253_n128, r253_n127, r253_n126,
         r253_n125, r253_n124, r253_n123, r253_n122, r253_n121, r253_n120,
         r253_n119, r253_n118, r253_n117, r253_n116, r253_n115, r253_n114,
         r253_n113, r253_n112, r253_n111, r253_n110, r253_n109, r253_n108,
         r253_n107, r253_n106, r253_n105, r253_n104, r253_n103, r253_n102,
         r253_n101, r253_n100, r253_n99, r253_n98, r253_n97, r253_n96,
         r253_n95, r253_n94, r253_n93, r253_n92, r253_n91, r253_n90, r253_n89,
         r253_n88, r253_n87, r253_n86, r253_n85, r253_n84, r253_n83, r253_n82,
         r253_n81, r253_n80, r253_n79, r253_n78, r253_n77, r253_n76, r253_n75,
         r253_n74, r253_n73, r253_n72, r253_n71, r253_n70, r253_n69, r253_n68,
         r253_n67, r253_n66, r253_n65, r253_n64, r253_n63, r253_n62, r253_n61,
         r253_n60, r253_n59, r253_n58, r253_n57, r253_n56, r253_n55, r253_n54,
         r253_n53, r253_n52, r253_n51, r253_n50, r253_n49, r253_n48, r253_n47,
         r253_n46, r253_n45, r253_n44, r253_n43, r253_n42, r253_n41, r253_n40,
         r253_n39, r253_n38, r253_n37, r253_n36, r253_n35, r253_n34, r253_n33,
         r253_n32, r253_n31, r253_n30, r253_n29, r253_n28, r253_n27, r253_n26,
         r253_n25, r253_n24, r253_n23, r253_n22, r253_n21, r253_n20, r253_n19,
         r253_n18, r253_n17, r253_n16, r253_n15, r253_n14, r253_n13, r253_n12,
         r253_n11, r253_n10, r253_n9, r253_n8, r253_n7, r253_n6, r253_n5,
         r253_n4, r253_n3, r253_n2, r253_n1, r1161_n15, r1161_n14, r1161_n13,
         r1161_n12, r1161_n11, r1161_n10, r1161_n9, r1161_n8, r1161_n7,
         r1161_n6, r1161_n5, r1161_n4, r1161_n3, r1161_n2, r1161_n1, r1158_n56,
         r1158_n55, r1158_n54, r1158_n53, r1158_n52, r1158_n51, r1158_n50,
         r1158_n49, r1158_n48, r1158_n47, r1158_n46, r1158_n45, r1158_n44,
         r1158_n43, r1158_n42, r1158_n41, r1158_n40, r1158_n39, r1158_n38,
         r1158_n37, r1158_n36, r1158_n35, r1158_n34, r1158_n33, r1158_n32,
         r1158_n31, r1158_n30, r1158_n29, r1158_n28, r1158_n27, r1158_n26,
         r1158_n25, r1158_n24, r1158_n23, r1158_n22, r1158_n21, r1158_n20,
         r1158_n19, r1158_n18, r1158_n17, r1158_n16, r1158_n15, r1158_n14,
         r1158_n13, r1158_n12, r1158_n11, r1158_n10, r1158_n9, r1158_n8,
         r1158_n7, r1158_n6, r1158_n5, r1158_n4, r1158_n3, r1158_n2, r1158_n1,
         r1160_n30, r1160_n29, r1160_n28, r1160_n27, r1160_n26, r1160_n25,
         r1160_n24, r1160_n23, r1160_n22, r1160_n21, r1160_n20, r1160_n19,
         r1160_n18, r1160_n17, r1160_n16, r1160_n15, r1160_n14, r1160_n13,
         r1160_n12, r1160_n11, r1160_n10, r1160_n9, r1160_n8, r1160_n7,
         r1160_n6, r1160_n5, r1160_n4, r1160_n3, r1160_n2, r1160_n1;
  wire   [31:0] rEIP;
  assign Datao[31] = 1'b0;

  FD2 RequestPending_reg ( .D(n3287), .CP(CLOCK), .CD(n567), .Q(n2217), .QN(
        n4451) );
  FD2 State_reg_2_ ( .D(n3286), .CP(CLOCK), .CD(n567), .Q(n2184), .QN(n4651)
         );
  FD2 State_reg_1_ ( .D(n3285), .CP(CLOCK), .CD(n567), .Q(n2150), .QN(n4667)
         );
  FD2 State_reg_0_ ( .D(n3284), .CP(CLOCK), .CD(n567), .Q(n4666), .QN(n2212)
         );
  FD2 DataWidth_reg_1_ ( .D(n3280), .CP(CLOCK), .CD(n567), .QN(n4656) );
  FD2 DataWidth_reg_0_ ( .D(n3281), .CP(CLOCK), .CD(n567), .QN(n4655) );
  FD2 StateBS16_reg ( .D(n3282), .CP(CLOCK), .CD(n567), .Q(n2214), .QN(n4665)
         );
  FD2 rEIP_reg_31_ ( .D(n3279), .CP(CLOCK), .CD(n567), .Q(rEIP[31]), .QN(n2154) );
  FD2 InstAddrPointer_reg_31_ ( .D(n3277), .CP(CLOCK), .CD(n567), .Q(n4657) );
  FD2 EBX_reg_1_ ( .D(n3194), .CP(CLOCK), .CD(n567), .QN(n4452) );
  FD2 rEIP_reg_1_ ( .D(n3267), .CP(CLOCK), .CD(n567), .Q(rEIP[1]), .QN(n2149)
         );
  FD2 InstAddrPointer_reg_1_ ( .D(n3002), .CP(CLOCK), .CD(n567), .Q(n4453) );
  FD2 InstQueueWr_Addr_reg_0_ ( .D(n3231), .CP(CLOCK), .CD(n567), .Q(n2169), 
        .QN(n4454) );
  FD2 InstQueueWr_Addr_reg_1_ ( .D(n3230), .CP(CLOCK), .CD(n567), .Q(n2146), 
        .QN(n4455) );
  FD2 InstQueueWr_Addr_reg_2_ ( .D(n3229), .CP(CLOCK), .CD(n567), .Q(n2147), 
        .QN(n4456) );
  FD2 InstQueueWr_Addr_reg_3_ ( .D(n3228), .CP(CLOCK), .CD(n567), .Q(n2171), 
        .QN(n4457) );
  FD2 State2_reg_0_ ( .D(n3275), .CP(CLOCK), .CD(n567), .Q(n2151), .QN(n4658)
         );
  FD2 State2_reg_1_ ( .D(n3273), .CP(CLOCK), .CD(n567), .QN(n4668) );
  FD2 State2_reg_3_ ( .D(n5488), .CP(CLOCK), .CD(n567), .Q(n2183), .QN(n4458)
         );
  FD2 State2_reg_2_ ( .D(n3274), .CP(CLOCK), .CD(n567), .Q(n2170), .QN(n4450)
         );
  FD2 PhyAddrPointer_reg_1_ ( .D(n2971), .CP(CLOCK), .CD(n567), .QN(n4459) );
  FD2 PhyAddrPointer_reg_0_ ( .D(n2972), .CP(CLOCK), .CD(n567), .QN(n4460) );
  FD2 rEIP_reg_0_ ( .D(n3268), .CP(CLOCK), .CD(n567), .Q(rEIP[0]), .QN(n2168)
         );
  FD2 InstAddrPointer_reg_0_ ( .D(n3003), .CP(CLOCK), .CD(n567), .Q(n4654) );
  FD2 InstQueueRd_Addr_reg_1_ ( .D(n3234), .CP(CLOCK), .CD(n567), .Q(n2167), 
        .QN(n4461) );
  FD2 CodeFetch_reg ( .D(n73), .CP(CLOCK), .CD(n567), .Q(n2216), .QN(n4652) );
  FD2 ReadRequest_reg ( .D(n3272), .CP(CLOCK), .CD(n567), .Q(n4354), .QN(n2215) );
  FD2 MemoryFetch_reg ( .D(n3270), .CP(CLOCK), .CD(n567), .QN(n4462) );
  FD2 Datao_reg_30_ ( .D(n2911), .CP(CLOCK), .CD(n567), .Q(Datao[30]), .QN(
        n5412) );
  FD2 Datao_reg_29_ ( .D(n2912), .CP(CLOCK), .CD(n567), .Q(Datao[29]), .QN(
        n5413) );
  FD2 Datao_reg_28_ ( .D(n2913), .CP(CLOCK), .CD(n567), .Q(Datao[28]), .QN(
        n5414) );
  FD2 Datao_reg_27_ ( .D(n2914), .CP(CLOCK), .CD(n567), .Q(Datao[27]), .QN(
        n5415) );
  FD2 Datao_reg_26_ ( .D(n2915), .CP(CLOCK), .CD(n567), .Q(Datao[26]), .QN(
        n5416) );
  FD2 Datao_reg_25_ ( .D(n2916), .CP(CLOCK), .CD(n567), .Q(Datao[25]), .QN(
        n5417) );
  FD2 Datao_reg_24_ ( .D(n2917), .CP(CLOCK), .CD(n567), .Q(Datao[24]), .QN(
        n5418) );
  FD2 Datao_reg_23_ ( .D(n2918), .CP(CLOCK), .CD(n567), .Q(Datao[23]), .QN(
        n5419) );
  FD2 Datao_reg_22_ ( .D(n2919), .CP(CLOCK), .CD(n567), .Q(Datao[22]), .QN(
        n5420) );
  FD2 Datao_reg_21_ ( .D(n2920), .CP(CLOCK), .CD(n567), .Q(Datao[21]), .QN(
        n5421) );
  FD2 Datao_reg_20_ ( .D(n2921), .CP(CLOCK), .CD(n567), .Q(Datao[20]), .QN(
        n5422) );
  FD2 Datao_reg_19_ ( .D(n2922), .CP(CLOCK), .CD(n567), .Q(Datao[19]), .QN(
        n5423) );
  FD2 Datao_reg_18_ ( .D(n2923), .CP(CLOCK), .CD(n567), .Q(Datao[18]), .QN(
        n5424) );
  FD2 Datao_reg_17_ ( .D(n2924), .CP(CLOCK), .CD(n567), .Q(Datao[17]), .QN(
        n5425) );
  FD2 Datao_reg_16_ ( .D(n2925), .CP(CLOCK), .CD(n567), .Q(Datao[16]), .QN(
        n5426) );
  FD2 EBX_reg_0_ ( .D(n3195), .CP(CLOCK), .CD(n567), .QN(n4463) );
  FD2 More_reg ( .D(n3004), .CP(CLOCK), .CD(n567), .QN(n4355) );
  FD2 Flush_reg ( .D(n22), .CP(CLOCK), .CD(n567), .QN(n4357) );
  FD2 EAX_reg_31_ ( .D(n3148), .CP(CLOCK), .CD(n567), .Q(n2197), .QN(n4464) );
  FD2 EAX_reg_0_ ( .D(n3210), .CP(CLOCK), .CD(n567), .Q(n4465) );
  FD2 Datao_reg_0_ ( .D(n2941), .CP(CLOCK), .CD(n567), .Q(Datao[0]), .QN(n5315) );
  FD2 lWord_reg_0_ ( .D(n3226), .CP(CLOCK), .CD(n567), .QN(n4466) );
  FD2 InstQueueRd_Addr_reg_3_ ( .D(n3276), .CP(CLOCK), .CD(n567), .Q(n2213), 
        .QN(n4467) );
  FD2 InstQueueRd_Addr_reg_0_ ( .D(n5489), .CP(CLOCK), .CD(n567), .Q(n2145), 
        .QN(n4468) );
  FD2 InstQueueRd_Addr_reg_2_ ( .D(n3233), .CP(CLOCK), .CD(n567), .Q(n2148), 
        .QN(n4653) );
  FD2 EAX_reg_1_ ( .D(n3209), .CP(CLOCK), .CD(n567), .Q(n4469) );
  FD2 Datao_reg_1_ ( .D(n2940), .CP(CLOCK), .CD(n567), .Q(Datao[1]), .QN(n5314) );
  FD2 lWord_reg_1_ ( .D(n3225), .CP(CLOCK), .CD(n567), .QN(n4470) );
  FD2 EBX_reg_2_ ( .D(n3193), .CP(CLOCK), .CD(n567), .QN(n4471) );
  FD2 rEIP_reg_2_ ( .D(n3266), .CP(CLOCK), .CD(n567), .Q(rEIP[2]), .QN(n2180)
         );
  FD2 PhyAddrPointer_reg_2_ ( .D(n2970), .CP(CLOCK), .CD(n567), .QN(n4472) );
  FD2 InstAddrPointer_reg_2_ ( .D(n3001), .CP(CLOCK), .CD(n567), .Q(n4473) );
  FD2 EAX_reg_2_ ( .D(n3208), .CP(CLOCK), .CD(n567), .Q(n4474) );
  FD2 Datao_reg_2_ ( .D(n2939), .CP(CLOCK), .CD(n567), .Q(Datao[2]), .QN(n5313) );
  FD2 lWord_reg_2_ ( .D(n3224), .CP(CLOCK), .CD(n567), .QN(n4475) );
  FD2 EBX_reg_3_ ( .D(n3192), .CP(CLOCK), .CD(n567), .QN(n4476) );
  FD2 rEIP_reg_3_ ( .D(n3265), .CP(CLOCK), .CD(n567), .Q(rEIP[3]), .QN(n2155)
         );
  FD2 PhyAddrPointer_reg_3_ ( .D(n2969), .CP(CLOCK), .CD(n567), .QN(n4477) );
  FD2 InstAddrPointer_reg_3_ ( .D(n3000), .CP(CLOCK), .CD(n567), .Q(n4478) );
  FD2 EAX_reg_3_ ( .D(n3207), .CP(CLOCK), .CD(n567), .Q(n4479) );
  FD2 Datao_reg_3_ ( .D(n2938), .CP(CLOCK), .CD(n567), .Q(Datao[3]), .QN(n5312) );
  FD2 lWord_reg_3_ ( .D(n3223), .CP(CLOCK), .CD(n567), .QN(n4480) );
  FD2 EBX_reg_4_ ( .D(n3191), .CP(CLOCK), .CD(n567), .QN(n4481) );
  FD2 rEIP_reg_4_ ( .D(n3264), .CP(CLOCK), .CD(n567), .Q(rEIP[4]), .QN(n2173)
         );
  FD2 PhyAddrPointer_reg_4_ ( .D(n2968), .CP(CLOCK), .CD(n567), .Q(n2185), 
        .QN(n4482) );
  FD2 InstAddrPointer_reg_4_ ( .D(n2999), .CP(CLOCK), .CD(n567), .Q(n4483) );
  FD2 EAX_reg_4_ ( .D(n3206), .CP(CLOCK), .CD(n567), .Q(n4484) );
  FD2 Datao_reg_4_ ( .D(n2937), .CP(CLOCK), .CD(n567), .Q(Datao[4]), .QN(n5311) );
  FD2 lWord_reg_4_ ( .D(n3222), .CP(CLOCK), .CD(n567), .QN(n4485) );
  FD2 EBX_reg_5_ ( .D(n3190), .CP(CLOCK), .CD(n567), .QN(n4486) );
  FD2 rEIP_reg_5_ ( .D(n3263), .CP(CLOCK), .CD(n567), .Q(rEIP[5]), .QN(n2153)
         );
  FD2 PhyAddrPointer_reg_5_ ( .D(n2967), .CP(CLOCK), .CD(n567), .Q(n2186), 
        .QN(n4487) );
  FD2 InstAddrPointer_reg_5_ ( .D(n2998), .CP(CLOCK), .CD(n567), .Q(n4488) );
  FD2 EAX_reg_5_ ( .D(n3205), .CP(CLOCK), .CD(n567), .Q(n4489) );
  FD2 Datao_reg_5_ ( .D(n2936), .CP(CLOCK), .CD(n567), .Q(Datao[5]), .QN(n5310) );
  FD2 lWord_reg_5_ ( .D(n3221), .CP(CLOCK), .CD(n567), .QN(n4490) );
  FD2 EBX_reg_6_ ( .D(n3189), .CP(CLOCK), .CD(n567), .Q(n2218), .QN(n4491) );
  FD2 rEIP_reg_6_ ( .D(n3262), .CP(CLOCK), .CD(n567), .Q(rEIP[6]), .QN(n2172)
         );
  FD2 PhyAddrPointer_reg_6_ ( .D(n2966), .CP(CLOCK), .CD(n567), .QN(n4492) );
  FD2 InstAddrPointer_reg_6_ ( .D(n2997), .CP(CLOCK), .CD(n567), .Q(n4493) );
  FD2 EAX_reg_6_ ( .D(n3204), .CP(CLOCK), .CD(n567), .Q(n4494) );
  FD2 Datao_reg_6_ ( .D(n2935), .CP(CLOCK), .CD(n567), .Q(Datao[6]), .QN(n5309) );
  FD2 lWord_reg_6_ ( .D(n3220), .CP(CLOCK), .CD(n567), .QN(n4495) );
  FD2 EBX_reg_7_ ( .D(n3188), .CP(CLOCK), .CD(n567), .Q(n2219), .QN(n4496) );
  FD2 rEIP_reg_7_ ( .D(n3261), .CP(CLOCK), .CD(n567), .Q(rEIP[7]), .QN(n2152)
         );
  FD2 PhyAddrPointer_reg_7_ ( .D(n2965), .CP(CLOCK), .CD(n567), .QN(n4497) );
  FD2 InstAddrPointer_reg_7_ ( .D(n2996), .CP(CLOCK), .CD(n567), .Q(n4498) );
  FD2 EAX_reg_7_ ( .D(n3203), .CP(CLOCK), .CD(n567), .Q(n4499) );
  FD2 Datao_reg_7_ ( .D(n2934), .CP(CLOCK), .CD(n567), .Q(Datao[7]), .QN(n5308) );
  FD2 lWord_reg_7_ ( .D(n3219), .CP(CLOCK), .CD(n567), .QN(n4500) );
  FD2 EBX_reg_8_ ( .D(n3187), .CP(CLOCK), .CD(n567), .Q(n2220), .QN(n4501) );
  FD2 rEIP_reg_8_ ( .D(n3260), .CP(CLOCK), .CD(n567), .Q(rEIP[8]), .QN(n2192)
         );
  FD2 PhyAddrPointer_reg_8_ ( .D(n2964), .CP(CLOCK), .CD(n567), .QN(n4502) );
  FD2 InstAddrPointer_reg_8_ ( .D(n2995), .CP(CLOCK), .CD(n567), .Q(n2196), 
        .QN(n4359) );
  FD2 EAX_reg_8_ ( .D(n3202), .CP(CLOCK), .CD(n567), .Q(n4503) );
  FD2 Datao_reg_8_ ( .D(n2933), .CP(CLOCK), .CD(n567), .Q(Datao[8]), .QN(n5307) );
  FD2 lWord_reg_8_ ( .D(n3218), .CP(CLOCK), .CD(n567), .QN(n4504) );
  FD2 EBX_reg_9_ ( .D(n3186), .CP(CLOCK), .CD(n567), .Q(n2221), .QN(n4505) );
  FD2 rEIP_reg_9_ ( .D(n3259), .CP(CLOCK), .CD(n567), .Q(rEIP[9]), .QN(n2163)
         );
  FD2 PhyAddrPointer_reg_9_ ( .D(n2963), .CP(CLOCK), .CD(n567), .QN(n4506) );
  FD2 InstAddrPointer_reg_9_ ( .D(n2994), .CP(CLOCK), .CD(n567), .Q(n2195), 
        .QN(n4358) );
  FD2 EAX_reg_9_ ( .D(n3201), .CP(CLOCK), .CD(n567), .Q(n4507) );
  FD2 Datao_reg_9_ ( .D(n2932), .CP(CLOCK), .CD(n567), .Q(Datao[9]), .QN(n5306) );
  FD2 lWord_reg_9_ ( .D(n3217), .CP(CLOCK), .CD(n567), .QN(n4508) );
  FD2 EBX_reg_10_ ( .D(n3185), .CP(CLOCK), .CD(n567), .Q(n2222), .QN(n4509) );
  FD2 rEIP_reg_10_ ( .D(n3258), .CP(CLOCK), .CD(n567), .Q(rEIP[10]), .QN(n2191) );
  FD2 PhyAddrPointer_reg_10_ ( .D(n2962), .CP(CLOCK), .CD(n567), .QN(n4510) );
  FD2 InstAddrPointer_reg_10_ ( .D(n2993), .CP(CLOCK), .CD(n567), .Q(n2211), 
        .QN(n4365) );
  FD2 EAX_reg_10_ ( .D(n3200), .CP(CLOCK), .CD(n567), .Q(n4511) );
  FD2 Datao_reg_10_ ( .D(n2931), .CP(CLOCK), .CD(n567), .Q(Datao[10]), .QN(
        n5305) );
  FD2 lWord_reg_10_ ( .D(n3216), .CP(CLOCK), .CD(n567), .QN(n4512) );
  FD2 EBX_reg_11_ ( .D(n3184), .CP(CLOCK), .CD(n567), .Q(n2223), .QN(n4513) );
  FD2 rEIP_reg_11_ ( .D(n3257), .CP(CLOCK), .CD(n567), .Q(rEIP[11]), .QN(n2166) );
  FD2 PhyAddrPointer_reg_11_ ( .D(n2961), .CP(CLOCK), .CD(n567), .QN(n4514) );
  FD2 InstAddrPointer_reg_11_ ( .D(n2992), .CP(CLOCK), .CD(n567), .Q(n2210), 
        .QN(n4364) );
  FD2 EAX_reg_11_ ( .D(n3199), .CP(CLOCK), .CD(n567), .Q(n4515) );
  FD2 Datao_reg_11_ ( .D(n2930), .CP(CLOCK), .CD(n567), .Q(Datao[11]), .QN(
        n5304) );
  FD2 lWord_reg_11_ ( .D(n3215), .CP(CLOCK), .CD(n567), .QN(n4516) );
  FD2 EBX_reg_12_ ( .D(n3183), .CP(CLOCK), .CD(n567), .Q(n2224), .QN(n4517) );
  FD2 rEIP_reg_12_ ( .D(n3256), .CP(CLOCK), .CD(n567), .Q(rEIP[12]), .QN(n2194) );
  FD2 PhyAddrPointer_reg_12_ ( .D(n2960), .CP(CLOCK), .CD(n567), .QN(n4518) );
  FD2 InstAddrPointer_reg_12_ ( .D(n2991), .CP(CLOCK), .CD(n567), .Q(n2209), 
        .QN(n4363) );
  FD2 EAX_reg_12_ ( .D(n3198), .CP(CLOCK), .CD(n567), .Q(n4519) );
  FD2 Datao_reg_12_ ( .D(n2929), .CP(CLOCK), .CD(n567), .Q(Datao[12]), .QN(
        n5303) );
  FD2 lWord_reg_12_ ( .D(n3214), .CP(CLOCK), .CD(n567), .QN(n4520) );
  FD2 EBX_reg_13_ ( .D(n3182), .CP(CLOCK), .CD(n567), .Q(n2225), .QN(n4521) );
  FD2 rEIP_reg_13_ ( .D(n3255), .CP(CLOCK), .CD(n567), .Q(rEIP[13]), .QN(n2165) );
  FD2 PhyAddrPointer_reg_13_ ( .D(n2959), .CP(CLOCK), .CD(n567), .QN(n4522) );
  FD2 InstAddrPointer_reg_13_ ( .D(n2990), .CP(CLOCK), .CD(n567), .Q(n2208), 
        .QN(n4362) );
  FD2 EAX_reg_13_ ( .D(n3197), .CP(CLOCK), .CD(n567), .Q(n4523) );
  FD2 Datao_reg_13_ ( .D(n2928), .CP(CLOCK), .CD(n567), .Q(Datao[13]), .QN(
        n5302) );
  FD2 lWord_reg_13_ ( .D(n3213), .CP(CLOCK), .CD(n567), .QN(n4524) );
  FD2 EBX_reg_14_ ( .D(n3181), .CP(CLOCK), .CD(n567), .Q(n2226), .QN(n4525) );
  FD2 rEIP_reg_14_ ( .D(n3254), .CP(CLOCK), .CD(n567), .Q(rEIP[14]), .QN(n2193) );
  FD2 PhyAddrPointer_reg_14_ ( .D(n2958), .CP(CLOCK), .CD(n567), .QN(n4526) );
  FD2 InstAddrPointer_reg_14_ ( .D(n2989), .CP(CLOCK), .CD(n567), .Q(n2207), 
        .QN(n4361) );
  FD2 EAX_reg_14_ ( .D(n3196), .CP(CLOCK), .CD(n567), .Q(n4527) );
  FD2 Datao_reg_14_ ( .D(n2927), .CP(CLOCK), .CD(n567), .Q(Datao[14]), .QN(
        n5301) );
  FD2 lWord_reg_14_ ( .D(n3212), .CP(CLOCK), .CD(n567), .QN(n4528) );
  FD2 EBX_reg_15_ ( .D(n3180), .CP(CLOCK), .CD(n567), .Q(n2227), .QN(n4529) );
  FD2 rEIP_reg_15_ ( .D(n3253), .CP(CLOCK), .CD(n567), .Q(rEIP[15]), .QN(n2164) );
  FD2 PhyAddrPointer_reg_15_ ( .D(n2957), .CP(CLOCK), .CD(n567), .QN(n4530) );
  FD2 InstAddrPointer_reg_15_ ( .D(n2988), .CP(CLOCK), .CD(n567), .Q(n2206), 
        .QN(n4360) );
  FD2 EAX_reg_15_ ( .D(n3227), .CP(CLOCK), .CD(n567), .Q(n4531) );
  FD2 Datao_reg_15_ ( .D(n2926), .CP(CLOCK), .CD(n567), .Q(Datao[15]), .QN(
        n5300) );
  FD2 lWord_reg_15_ ( .D(n3211), .CP(CLOCK), .CD(n567), .QN(n4532) );
  FD2 EAX_reg_16_ ( .D(n3163), .CP(CLOCK), .CD(n567), .Q(n4533) );
  FD2 EBX_reg_16_ ( .D(n3179), .CP(CLOCK), .CD(n567), .Q(n2190), .QN(n4534) );
  FD2 rEIP_reg_16_ ( .D(n3252), .CP(CLOCK), .CD(n567), .Q(rEIP[16]), .QN(n2182) );
  FD2 PhyAddrPointer_reg_16_ ( .D(n2956), .CP(CLOCK), .CD(n567), .QN(n4535) );
  FD2 InstAddrPointer_reg_16_ ( .D(n2987), .CP(CLOCK), .CD(n567), .Q(n4536) );
  FD2 EAX_reg_17_ ( .D(n3162), .CP(CLOCK), .CD(n567), .Q(n4537) );
  FD2 EBX_reg_17_ ( .D(n3178), .CP(CLOCK), .CD(n567), .Q(n2189), .QN(n4538) );
  FD2 rEIP_reg_17_ ( .D(n3251), .CP(CLOCK), .CD(n567), .Q(rEIP[17]), .QN(n2162) );
  FD2 PhyAddrPointer_reg_17_ ( .D(n2955), .CP(CLOCK), .CD(n567), .QN(n4539) );
  FD2 InstAddrPointer_reg_17_ ( .D(n2986), .CP(CLOCK), .CD(n567), .Q(n4540) );
  FD2 EAX_reg_18_ ( .D(n3161), .CP(CLOCK), .CD(n567), .Q(n4541) );
  FD2 EBX_reg_18_ ( .D(n3177), .CP(CLOCK), .CD(n567), .Q(n2188), .QN(n4542) );
  FD2 rEIP_reg_18_ ( .D(n3250), .CP(CLOCK), .CD(n567), .Q(rEIP[18]), .QN(n2181) );
  FD2 PhyAddrPointer_reg_18_ ( .D(n2954), .CP(CLOCK), .CD(n567), .QN(n4543) );
  FD2 InstAddrPointer_reg_18_ ( .D(n2985), .CP(CLOCK), .CD(n567), .Q(n4544) );
  FD2 EAX_reg_19_ ( .D(n3160), .CP(CLOCK), .CD(n567), .Q(n4545) );
  FD2 EBX_reg_19_ ( .D(n3176), .CP(CLOCK), .CD(n567), .Q(n2187), .QN(n4546) );
  FD2 rEIP_reg_19_ ( .D(n3249), .CP(CLOCK), .CD(n567), .Q(rEIP[19]), .QN(n2161) );
  FD2 PhyAddrPointer_reg_19_ ( .D(n2953), .CP(CLOCK), .CD(n567), .QN(n4547) );
  FD2 InstAddrPointer_reg_19_ ( .D(n2984), .CP(CLOCK), .CD(n567), .Q(n4548) );
  FD2 EAX_reg_20_ ( .D(n3159), .CP(CLOCK), .CD(n567), .Q(n4549) );
  FD2 EBX_reg_20_ ( .D(n3175), .CP(CLOCK), .CD(n567), .QN(n4550) );
  FD2 rEIP_reg_20_ ( .D(n3248), .CP(CLOCK), .CD(n567), .Q(rEIP[20]), .QN(n2179) );
  FD2 PhyAddrPointer_reg_20_ ( .D(n2952), .CP(CLOCK), .CD(n567), .QN(n4551) );
  FD2 InstAddrPointer_reg_20_ ( .D(n2983), .CP(CLOCK), .CD(n567), .Q(n4552) );
  FD2 EAX_reg_21_ ( .D(n3158), .CP(CLOCK), .CD(n567), .Q(n4553) );
  FD2 EBX_reg_21_ ( .D(n3174), .CP(CLOCK), .CD(n567), .QN(n4554) );
  FD2 rEIP_reg_21_ ( .D(n3247), .CP(CLOCK), .CD(n567), .Q(rEIP[21]), .QN(n2160) );
  FD2 PhyAddrPointer_reg_21_ ( .D(n2951), .CP(CLOCK), .CD(n567), .QN(n4555) );
  FD2 InstAddrPointer_reg_21_ ( .D(n2982), .CP(CLOCK), .CD(n567), .Q(n4556) );
  FD2 EAX_reg_22_ ( .D(n3157), .CP(CLOCK), .CD(n567), .Q(n4557) );
  FD2 EBX_reg_22_ ( .D(n3173), .CP(CLOCK), .CD(n567), .QN(n4558) );
  FD2 rEIP_reg_22_ ( .D(n3246), .CP(CLOCK), .CD(n567), .Q(rEIP[22]), .QN(n2178) );
  FD2 PhyAddrPointer_reg_22_ ( .D(n2950), .CP(CLOCK), .CD(n567), .QN(n4559) );
  FD2 InstAddrPointer_reg_22_ ( .D(n2981), .CP(CLOCK), .CD(n567), .Q(n4560) );
  FD2 EAX_reg_23_ ( .D(n3156), .CP(CLOCK), .CD(n567), .Q(n2205), .QN(n4561) );
  FD2 EBX_reg_23_ ( .D(n3172), .CP(CLOCK), .CD(n567), .QN(n4562) );
  FD2 rEIP_reg_23_ ( .D(n3245), .CP(CLOCK), .CD(n567), .Q(rEIP[23]), .QN(n2159) );
  FD2 PhyAddrPointer_reg_23_ ( .D(n2949), .CP(CLOCK), .CD(n567), .QN(n4563) );
  FD2 InstAddrPointer_reg_23_ ( .D(n2980), .CP(CLOCK), .CD(n567), .Q(n4564) );
  FD2 EAX_reg_24_ ( .D(n3155), .CP(CLOCK), .CD(n567), .Q(n2204), .QN(n4565) );
  FD2 EBX_reg_24_ ( .D(n3171), .CP(CLOCK), .CD(n567), .QN(n4566) );
  FD2 rEIP_reg_24_ ( .D(n3244), .CP(CLOCK), .CD(n567), .Q(rEIP[24]), .QN(n2177) );
  FD2 PhyAddrPointer_reg_24_ ( .D(n2948), .CP(CLOCK), .CD(n567), .QN(n4567) );
  FD2 InstAddrPointer_reg_24_ ( .D(n2979), .CP(CLOCK), .CD(n567), .Q(n4568) );
  FD2 EAX_reg_25_ ( .D(n3154), .CP(CLOCK), .CD(n567), .Q(n2203), .QN(n4569) );
  FD2 EBX_reg_25_ ( .D(n3170), .CP(CLOCK), .CD(n567), .QN(n4570) );
  FD2 rEIP_reg_25_ ( .D(n3243), .CP(CLOCK), .CD(n567), .Q(rEIP[25]), .QN(n2158) );
  FD2 PhyAddrPointer_reg_25_ ( .D(n2947), .CP(CLOCK), .CD(n567), .QN(n4571) );
  FD2 InstAddrPointer_reg_25_ ( .D(n2978), .CP(CLOCK), .CD(n567), .Q(n4572) );
  FD2 EAX_reg_26_ ( .D(n3153), .CP(CLOCK), .CD(n567), .Q(n2202), .QN(n4573) );
  FD2 EBX_reg_26_ ( .D(n3169), .CP(CLOCK), .CD(n567), .QN(n4574) );
  FD2 rEIP_reg_26_ ( .D(n3242), .CP(CLOCK), .CD(n567), .Q(rEIP[26]), .QN(n2176) );
  FD2 PhyAddrPointer_reg_26_ ( .D(n2946), .CP(CLOCK), .CD(n567), .QN(n4575) );
  FD2 InstAddrPointer_reg_26_ ( .D(n2977), .CP(CLOCK), .CD(n567), .Q(n4576) );
  FD2 EAX_reg_27_ ( .D(n3152), .CP(CLOCK), .CD(n567), .Q(n2201), .QN(n4577) );
  FD2 EBX_reg_27_ ( .D(n3168), .CP(CLOCK), .CD(n567), .QN(n4578) );
  FD2 rEIP_reg_27_ ( .D(n3241), .CP(CLOCK), .CD(n567), .Q(rEIP[27]), .QN(n2157) );
  FD2 PhyAddrPointer_reg_27_ ( .D(n2945), .CP(CLOCK), .CD(n567), .QN(n4579) );
  FD2 InstAddrPointer_reg_27_ ( .D(n2976), .CP(CLOCK), .CD(n567), .Q(n4580) );
  FD2 EAX_reg_28_ ( .D(n3151), .CP(CLOCK), .CD(n567), .Q(n2200), .QN(n4581) );
  FD2 EBX_reg_28_ ( .D(n3167), .CP(CLOCK), .CD(n567), .QN(n4582) );
  FD2 rEIP_reg_28_ ( .D(n3240), .CP(CLOCK), .CD(n567), .Q(rEIP[28]), .QN(n2175) );
  FD2 PhyAddrPointer_reg_28_ ( .D(n2944), .CP(CLOCK), .CD(n567), .QN(n4583) );
  FD2 InstAddrPointer_reg_28_ ( .D(n2975), .CP(CLOCK), .CD(n567), .Q(n4584) );
  FD2 EAX_reg_29_ ( .D(n3150), .CP(CLOCK), .CD(n567), .Q(n2199), .QN(n4585) );
  FD2 EBX_reg_29_ ( .D(n3166), .CP(CLOCK), .CD(n567), .QN(n4586) );
  FD2 rEIP_reg_29_ ( .D(n3239), .CP(CLOCK), .CD(n567), .Q(rEIP[29]), .QN(n2156) );
  FD2 PhyAddrPointer_reg_29_ ( .D(n2943), .CP(CLOCK), .CD(n567), .QN(n4587) );
  FD2 InstAddrPointer_reg_29_ ( .D(n2974), .CP(CLOCK), .CD(n567), .Q(n4588) );
  FD2 EAX_reg_30_ ( .D(n3149), .CP(CLOCK), .CD(n567), .Q(n2198), .QN(n4589) );
  FD2 uWord_reg_0_ ( .D(n3019), .CP(CLOCK), .CD(n567), .QN(n4590) );
  FD2 InstQueue_reg_15__0_ ( .D(n3027), .CP(CLOCK), .CD(n567), .Q(n4409) );
  FD2 InstQueue_reg_14__0_ ( .D(n3035), .CP(CLOCK), .CD(n567), .Q(n4406) );
  FD2 InstQueue_reg_13__0_ ( .D(n3043), .CP(CLOCK), .CD(n567), .Q(n4415) );
  FD2 InstQueue_reg_12__0_ ( .D(n3051), .CP(CLOCK), .CD(n567), .Q(n4414) );
  FD2 InstQueue_reg_11__0_ ( .D(n3059), .CP(CLOCK), .CD(n567), .Q(n4411) );
  FD2 InstQueue_reg_10__0_ ( .D(n3067), .CP(CLOCK), .CD(n567), .Q(n4408) );
  FD2 InstQueue_reg_9__0_ ( .D(n3075), .CP(CLOCK), .CD(n567), .Q(n4417), .QN(
        n2237) );
  FD2 InstQueue_reg_8__0_ ( .D(n3083), .CP(CLOCK), .CD(n567), .Q(n4591) );
  FD2 InstQueue_reg_7__0_ ( .D(n3091), .CP(CLOCK), .CD(n567), .Q(n4592) );
  FD2 InstQueue_reg_6__0_ ( .D(n3099), .CP(CLOCK), .CD(n567), .Q(n4593) );
  FD2 InstQueue_reg_5__0_ ( .D(n3107), .CP(CLOCK), .CD(n567), .Q(n4594) );
  FD2 InstQueue_reg_4__0_ ( .D(n3115), .CP(CLOCK), .CD(n567), .Q(n4412) );
  FD2 InstQueue_reg_3__0_ ( .D(n3123), .CP(CLOCK), .CD(n567), .Q(n4410) );
  FD2 InstQueue_reg_2__0_ ( .D(n3131), .CP(CLOCK), .CD(n567), .Q(n4407) );
  FD2 InstQueue_reg_1__0_ ( .D(n3139), .CP(CLOCK), .CD(n567), .Q(n4416) );
  FD2 InstQueue_reg_0__0_ ( .D(n3147), .CP(CLOCK), .CD(n567), .Q(n4413) );
  FD2 uWord_reg_1_ ( .D(n3018), .CP(CLOCK), .CD(n567), .QN(n4595) );
  FD2 InstQueue_reg_15__1_ ( .D(n3026), .CP(CLOCK), .CD(n567), .Q(n4421) );
  FD2 InstQueue_reg_14__1_ ( .D(n3034), .CP(CLOCK), .CD(n567), .Q(n4418) );
  FD2 InstQueue_reg_13__1_ ( .D(n3042), .CP(CLOCK), .CD(n567), .Q(n4427) );
  FD2 InstQueue_reg_12__1_ ( .D(n3050), .CP(CLOCK), .CD(n567), .Q(n4426) );
  FD2 InstQueue_reg_11__1_ ( .D(n3058), .CP(CLOCK), .CD(n567), .Q(n4423), .QN(
        n2230) );
  FD2 InstQueue_reg_10__1_ ( .D(n3066), .CP(CLOCK), .CD(n567), .Q(n4420) );
  FD2 InstQueue_reg_9__1_ ( .D(n3074), .CP(CLOCK), .CD(n567), .Q(n4429) );
  FD2 InstQueue_reg_8__1_ ( .D(n3082), .CP(CLOCK), .CD(n567), .Q(n4596) );
  FD2 InstQueue_reg_7__1_ ( .D(n3090), .CP(CLOCK), .CD(n567), .Q(n4597) );
  FD2 InstQueue_reg_6__1_ ( .D(n3098), .CP(CLOCK), .CD(n567), .Q(n4598) );
  FD2 InstQueue_reg_5__1_ ( .D(n3106), .CP(CLOCK), .CD(n567), .Q(n4599) );
  FD2 InstQueue_reg_4__1_ ( .D(n3114), .CP(CLOCK), .CD(n567), .Q(n4424) );
  FD2 InstQueue_reg_3__1_ ( .D(n3122), .CP(CLOCK), .CD(n567), .Q(n4422) );
  FD2 InstQueue_reg_2__1_ ( .D(n3130), .CP(CLOCK), .CD(n567), .Q(n4419) );
  FD2 InstQueue_reg_1__1_ ( .D(n3138), .CP(CLOCK), .CD(n567), .Q(n4428) );
  FD2 InstQueue_reg_0__1_ ( .D(n3146), .CP(CLOCK), .CD(n567), .Q(n4425) );
  FD2 uWord_reg_2_ ( .D(n3017), .CP(CLOCK), .CD(n567), .QN(n4600) );
  FD2 InstQueue_reg_15__2_ ( .D(n3025), .CP(CLOCK), .CD(n567), .Q(n4399) );
  FD2 InstQueue_reg_14__2_ ( .D(n3033), .CP(CLOCK), .CD(n567), .Q(n4396) );
  FD2 InstQueue_reg_13__2_ ( .D(n3041), .CP(CLOCK), .CD(n567), .Q(n4404) );
  FD2 InstQueue_reg_12__2_ ( .D(n3049), .CP(CLOCK), .CD(n567), .Q(n4403) );
  FD2 InstQueue_reg_11__2_ ( .D(n3057), .CP(CLOCK), .CD(n567), .Q(n4401), .QN(
        n2229) );
  FD2 InstQueue_reg_10__2_ ( .D(n3065), .CP(CLOCK), .CD(n567), .Q(n4398) );
  FD2 InstQueue_reg_9__2_ ( .D(n3073), .CP(CLOCK), .CD(n567), .Q(n4601) );
  FD2 InstQueue_reg_8__2_ ( .D(n3081), .CP(CLOCK), .CD(n567), .Q(n4602) );
  FD2 InstQueue_reg_7__2_ ( .D(n3089), .CP(CLOCK), .CD(n567), .Q(n4603) );
  FD2 InstQueue_reg_6__2_ ( .D(n3097), .CP(CLOCK), .CD(n567), .Q(n4604) );
  FD2 InstQueue_reg_5__2_ ( .D(n3105), .CP(CLOCK), .CD(n567), .Q(n4605) );
  FD2 InstQueue_reg_4__2_ ( .D(n3113), .CP(CLOCK), .CD(n567), .Q(n4402) );
  FD2 InstQueue_reg_3__2_ ( .D(n3121), .CP(CLOCK), .CD(n567), .Q(n4400) );
  FD2 InstQueue_reg_2__2_ ( .D(n3129), .CP(CLOCK), .CD(n567), .Q(n4397) );
  FD2 InstQueue_reg_1__2_ ( .D(n3137), .CP(CLOCK), .CD(n567), .Q(n4405) );
  FD2 InstQueue_reg_0__2_ ( .D(n3145), .CP(CLOCK), .CD(n567), .Q(n4664), .QN(
        n2236) );
  FD2 uWord_reg_3_ ( .D(n3016), .CP(CLOCK), .CD(n567), .QN(n4606) );
  FD2 InstQueue_reg_15__3_ ( .D(n3024), .CP(CLOCK), .CD(n567), .Q(n4432) );
  FD2 InstQueue_reg_14__3_ ( .D(n3032), .CP(CLOCK), .CD(n567), .Q(n4430) );
  FD2 InstQueue_reg_13__3_ ( .D(n3040), .CP(CLOCK), .CD(n567), .Q(n4437) );
  FD2 InstQueue_reg_12__3_ ( .D(n3048), .CP(CLOCK), .CD(n567), .Q(n4436) );
  FD2 InstQueue_reg_11__3_ ( .D(n3056), .CP(CLOCK), .CD(n567), .Q(n4434) );
  FD2 InstQueue_reg_10__3_ ( .D(n3064), .CP(CLOCK), .CD(n567), .Q(n4607) );
  FD2 InstQueue_reg_9__3_ ( .D(n3072), .CP(CLOCK), .CD(n567), .Q(n4439) );
  FD2 InstQueue_reg_8__3_ ( .D(n3080), .CP(CLOCK), .CD(n567), .Q(n4608), .QN(
        n2241) );
  FD2 InstQueue_reg_7__3_ ( .D(n3088), .CP(CLOCK), .CD(n567), .Q(n4609) );
  FD2 InstQueue_reg_6__3_ ( .D(n3096), .CP(CLOCK), .CD(n567), .Q(n4610) );
  FD2 InstQueue_reg_5__3_ ( .D(n3104), .CP(CLOCK), .CD(n567), .Q(n4611) );
  FD2 InstQueue_reg_4__3_ ( .D(n3112), .CP(CLOCK), .CD(n567), .Q(n4435) );
  FD2 InstQueue_reg_3__3_ ( .D(n3120), .CP(CLOCK), .CD(n567), .Q(n4433) );
  FD2 InstQueue_reg_2__3_ ( .D(n3128), .CP(CLOCK), .CD(n567), .Q(n4431) );
  FD2 InstQueue_reg_1__3_ ( .D(n3136), .CP(CLOCK), .CD(n567), .Q(n4438) );
  FD2 InstQueue_reg_0__3_ ( .D(n3144), .CP(CLOCK), .CD(n567), .Q(n4663), .QN(
        n2235) );
  FD2 uWord_reg_4_ ( .D(n3015), .CP(CLOCK), .CD(n567), .QN(n4612) );
  FD2 InstQueue_reg_15__4_ ( .D(n3023), .CP(CLOCK), .CD(n567), .Q(n4442) );
  FD2 InstQueue_reg_14__4_ ( .D(n3031), .CP(CLOCK), .CD(n567), .Q(n4440) );
  FD2 InstQueue_reg_13__4_ ( .D(n3039), .CP(CLOCK), .CD(n567), .Q(n4447) );
  FD2 InstQueue_reg_12__4_ ( .D(n3047), .CP(CLOCK), .CD(n567), .Q(n4446) );
  FD2 InstQueue_reg_11__4_ ( .D(n3055), .CP(CLOCK), .CD(n567), .Q(n4444) );
  FD2 InstQueue_reg_10__4_ ( .D(n3063), .CP(CLOCK), .CD(n567), .Q(n4613) );
  FD2 InstQueue_reg_9__4_ ( .D(n3071), .CP(CLOCK), .CD(n567), .Q(n4449) );
  FD2 InstQueue_reg_8__4_ ( .D(n3079), .CP(CLOCK), .CD(n567), .Q(n4614), .QN(
        n2240) );
  FD2 InstQueue_reg_7__4_ ( .D(n3087), .CP(CLOCK), .CD(n567), .Q(n4615) );
  FD2 InstQueue_reg_6__4_ ( .D(n3095), .CP(CLOCK), .CD(n567), .Q(n4616) );
  FD2 InstQueue_reg_5__4_ ( .D(n3103), .CP(CLOCK), .CD(n567), .Q(n4617) );
  FD2 InstQueue_reg_4__4_ ( .D(n3111), .CP(CLOCK), .CD(n567), .Q(n4445) );
  FD2 InstQueue_reg_3__4_ ( .D(n3119), .CP(CLOCK), .CD(n567), .Q(n4443) );
  FD2 InstQueue_reg_2__4_ ( .D(n3127), .CP(CLOCK), .CD(n567), .Q(n4441) );
  FD2 InstQueue_reg_1__4_ ( .D(n3135), .CP(CLOCK), .CD(n567), .Q(n4448) );
  FD2 InstQueue_reg_0__4_ ( .D(n3143), .CP(CLOCK), .CD(n567), .Q(n4662), .QN(
        n2234) );
  FD2 uWord_reg_5_ ( .D(n3014), .CP(CLOCK), .CD(n567), .QN(n4618) );
  FD2 InstQueue_reg_15__5_ ( .D(n3022), .CP(CLOCK), .CD(n567), .Q(n4368) );
  FD2 InstQueue_reg_14__5_ ( .D(n3030), .CP(CLOCK), .CD(n567), .Q(n4366) );
  FD2 InstQueue_reg_13__5_ ( .D(n3038), .CP(CLOCK), .CD(n567), .Q(n4373) );
  FD2 InstQueue_reg_12__5_ ( .D(n3046), .CP(CLOCK), .CD(n567), .Q(n4372) );
  FD2 InstQueue_reg_11__5_ ( .D(n3054), .CP(CLOCK), .CD(n567), .Q(n4370) );
  FD2 InstQueue_reg_10__5_ ( .D(n3062), .CP(CLOCK), .CD(n567), .Q(n4619) );
  FD2 InstQueue_reg_9__5_ ( .D(n3070), .CP(CLOCK), .CD(n567), .Q(n4375) );
  FD2 InstQueue_reg_8__5_ ( .D(n3078), .CP(CLOCK), .CD(n567), .Q(n4620), .QN(
        n2239) );
  FD2 InstQueue_reg_7__5_ ( .D(n3086), .CP(CLOCK), .CD(n567), .Q(n4621) );
  FD2 InstQueue_reg_6__5_ ( .D(n3094), .CP(CLOCK), .CD(n567), .Q(n4622) );
  FD2 InstQueue_reg_5__5_ ( .D(n3102), .CP(CLOCK), .CD(n567), .Q(n4623) );
  FD2 InstQueue_reg_4__5_ ( .D(n3110), .CP(CLOCK), .CD(n567), .Q(n4371) );
  FD2 InstQueue_reg_3__5_ ( .D(n3118), .CP(CLOCK), .CD(n567), .Q(n4369) );
  FD2 InstQueue_reg_2__5_ ( .D(n3126), .CP(CLOCK), .CD(n567), .Q(n4367) );
  FD2 InstQueue_reg_1__5_ ( .D(n3134), .CP(CLOCK), .CD(n567), .Q(n4374) );
  FD2 InstQueue_reg_0__5_ ( .D(n3142), .CP(CLOCK), .CD(n567), .Q(n4661), .QN(
        n2233) );
  FD2 uWord_reg_6_ ( .D(n3013), .CP(CLOCK), .CD(n567), .QN(n4624) );
  FD2 InstQueue_reg_15__6_ ( .D(n3021), .CP(CLOCK), .CD(n567), .Q(n4389) );
  FD2 InstQueue_reg_14__6_ ( .D(n3029), .CP(CLOCK), .CD(n567), .Q(n4387) );
  FD2 InstQueue_reg_13__6_ ( .D(n3037), .CP(CLOCK), .CD(n567), .Q(n4394) );
  FD2 InstQueue_reg_12__6_ ( .D(n3045), .CP(CLOCK), .CD(n567), .Q(n4393) );
  FD2 InstQueue_reg_11__6_ ( .D(n3053), .CP(CLOCK), .CD(n567), .Q(n4391) );
  FD2 InstQueue_reg_10__6_ ( .D(n3061), .CP(CLOCK), .CD(n567), .Q(n4625) );
  FD2 InstQueue_reg_9__6_ ( .D(n3069), .CP(CLOCK), .CD(n567), .Q(n4626) );
  FD2 InstQueue_reg_8__6_ ( .D(n3077), .CP(CLOCK), .CD(n567), .Q(n4627), .QN(
        n2238) );
  FD2 InstQueue_reg_7__6_ ( .D(n3085), .CP(CLOCK), .CD(n567), .Q(n4628) );
  FD2 InstQueue_reg_6__6_ ( .D(n3093), .CP(CLOCK), .CD(n567), .Q(n4629) );
  FD2 InstQueue_reg_5__6_ ( .D(n3101), .CP(CLOCK), .CD(n567), .Q(n4630) );
  FD2 InstQueue_reg_4__6_ ( .D(n3109), .CP(CLOCK), .CD(n567), .Q(n4392) );
  FD2 InstQueue_reg_3__6_ ( .D(n3117), .CP(CLOCK), .CD(n567), .Q(n4390) );
  FD2 InstQueue_reg_2__6_ ( .D(n3125), .CP(CLOCK), .CD(n567), .Q(n4388) );
  FD2 InstQueue_reg_1__6_ ( .D(n3133), .CP(CLOCK), .CD(n567), .Q(n4395) );
  FD2 InstQueue_reg_0__6_ ( .D(n3141), .CP(CLOCK), .CD(n567), .Q(n4660), .QN(
        n2232) );
  FD2 uWord_reg_7_ ( .D(n3012), .CP(CLOCK), .CD(n567), .QN(n4631) );
  FD2 InstQueue_reg_15__7_ ( .D(n35), .CP(CLOCK), .CD(n567), .Q(n4379) );
  FD2 InstQueue_reg_14__7_ ( .D(n3028), .CP(CLOCK), .CD(n567), .Q(n4376) );
  FD2 InstQueue_reg_13__7_ ( .D(n3036), .CP(CLOCK), .CD(n567), .Q(n4384) );
  FD2 InstQueue_reg_12__7_ ( .D(n3044), .CP(CLOCK), .CD(n567), .Q(n4383) );
  FD2 InstQueue_reg_11__7_ ( .D(n3052), .CP(CLOCK), .CD(n567), .Q(n4381), .QN(
        n2228) );
  FD2 InstQueue_reg_10__7_ ( .D(n3060), .CP(CLOCK), .CD(n567), .Q(n4378) );
  FD2 InstQueue_reg_9__7_ ( .D(n3068), .CP(CLOCK), .CD(n567), .Q(n4386) );
  FD2 InstQueue_reg_8__7_ ( .D(n3076), .CP(CLOCK), .CD(n567), .Q(n4632) );
  FD2 InstQueue_reg_7__7_ ( .D(n3084), .CP(CLOCK), .CD(n567), .Q(n4633) );
  FD2 InstQueue_reg_6__7_ ( .D(n3092), .CP(CLOCK), .CD(n567), .Q(n4634) );
  FD2 InstQueue_reg_5__7_ ( .D(n3100), .CP(CLOCK), .CD(n567), .Q(n4635) );
  FD2 InstQueue_reg_4__7_ ( .D(n3108), .CP(CLOCK), .CD(n567), .Q(n4382) );
  FD2 InstQueue_reg_3__7_ ( .D(n3116), .CP(CLOCK), .CD(n567), .Q(n4380) );
  FD2 InstQueue_reg_2__7_ ( .D(n3124), .CP(CLOCK), .CD(n567), .Q(n4377) );
  FD2 InstQueue_reg_1__7_ ( .D(n3132), .CP(CLOCK), .CD(n567), .Q(n4385) );
  FD2 InstQueue_reg_0__7_ ( .D(n3140), .CP(CLOCK), .CD(n567), .Q(n4659), .QN(
        n2231) );
  FD2 uWord_reg_8_ ( .D(n3011), .CP(CLOCK), .CD(n567), .QN(n4636) );
  FD2 uWord_reg_9_ ( .D(n3010), .CP(CLOCK), .CD(n567), .QN(n4637) );
  FD2 uWord_reg_10_ ( .D(n3009), .CP(CLOCK), .CD(n567), .QN(n4638) );
  FD2 uWord_reg_11_ ( .D(n3008), .CP(CLOCK), .CD(n567), .QN(n4639) );
  FD2 uWord_reg_12_ ( .D(n3007), .CP(CLOCK), .CD(n567), .QN(n4640) );
  FD2 uWord_reg_13_ ( .D(n3006), .CP(CLOCK), .CD(n567), .QN(n4641) );
  FD2 uWord_reg_14_ ( .D(n3005), .CP(CLOCK), .CD(n567), .QN(n4642) );
  FD2 EBX_reg_30_ ( .D(n3165), .CP(CLOCK), .CD(n567), .QN(n4643) );
  FD2 rEIP_reg_30_ ( .D(n3238), .CP(CLOCK), .CD(n567), .Q(rEIP[30]), .QN(n2174) );
  FD2 PhyAddrPointer_reg_30_ ( .D(n2942), .CP(CLOCK), .CD(n567), .QN(n4644) );
  FD2 InstAddrPointer_reg_30_ ( .D(n2973), .CP(CLOCK), .CD(n567), .Q(n4645) );
  FD2 EBX_reg_31_ ( .D(n3164), .CP(CLOCK), .CD(n567), .QN(n4646) );
  FD2 PhyAddrPointer_reg_31_ ( .D(n3278), .CP(CLOCK), .CD(n567), .QN(n4647) );
  FD2 W_R_n_reg ( .D(n3271), .CP(CLOCK), .CD(n567), .Q(W_R_n), .QN(n5430) );
  FD2 M_IO_n_reg ( .D(n3269), .CP(CLOCK), .CD(n567), .Q(M_IO_n), .QN(n5429) );
  FD2 D_C_n_reg ( .D(n3236), .CP(CLOCK), .CD(n567), .Q(D_C_n) );
  FD2 ADS_n_reg ( .D(n3283), .CP(CLOCK), .CD(n567), .Q(ADS_n), .QN(n5397) );
  FD2 Address_reg_0_ ( .D(n5521), .CP(CLOCK), .CD(n567), .Q(Address[0]) );
  FD2 Address_reg_1_ ( .D(n5492), .CP(CLOCK), .CD(n567), .Q(Address[1]) );
  FD2 Address_reg_2_ ( .D(n5519), .CP(CLOCK), .CD(n567), .Q(Address[2]) );
  FD2 Address_reg_3_ ( .D(n5520), .CP(CLOCK), .CD(n567), .Q(Address[3]) );
  FD2 Address_reg_4_ ( .D(n5517), .CP(CLOCK), .CD(n567), .Q(Address[4]) );
  FD2 Address_reg_5_ ( .D(n5518), .CP(CLOCK), .CD(n567), .Q(Address[5]) );
  FD2 Address_reg_6_ ( .D(n5515), .CP(CLOCK), .CD(n567), .Q(Address[6]) );
  FD2 Address_reg_7_ ( .D(n5516), .CP(CLOCK), .CD(n567), .Q(Address[7]) );
  FD2 Address_reg_8_ ( .D(n5513), .CP(CLOCK), .CD(n567), .Q(Address[8]) );
  FD2 Address_reg_9_ ( .D(n5514), .CP(CLOCK), .CD(n567), .Q(Address[9]) );
  FD2 Address_reg_10_ ( .D(n5493), .CP(CLOCK), .CD(n567), .Q(Address[10]) );
  FD2 Address_reg_11_ ( .D(n5494), .CP(CLOCK), .CD(n567), .Q(Address[11]) );
  FD2 Address_reg_12_ ( .D(n5495), .CP(CLOCK), .CD(n567), .Q(Address[12]) );
  FD2 Address_reg_13_ ( .D(n5496), .CP(CLOCK), .CD(n567), .Q(Address[13]) );
  FD2 Address_reg_14_ ( .D(n5497), .CP(CLOCK), .CD(n567), .Q(Address[14]) );
  FD2 Address_reg_15_ ( .D(n5498), .CP(CLOCK), .CD(n567), .Q(Address[15]) );
  FD2 Address_reg_16_ ( .D(n5499), .CP(CLOCK), .CD(n567), .Q(Address[16]) );
  FD2 Address_reg_17_ ( .D(n5500), .CP(CLOCK), .CD(n567), .Q(Address[17]) );
  FD2 Address_reg_18_ ( .D(n5501), .CP(CLOCK), .CD(n567), .Q(Address[18]) );
  FD2 Address_reg_19_ ( .D(n5502), .CP(CLOCK), .CD(n567), .Q(Address[19]) );
  FD2 Address_reg_20_ ( .D(n5503), .CP(CLOCK), .CD(n567), .Q(Address[20]) );
  FD2 Address_reg_21_ ( .D(n5504), .CP(CLOCK), .CD(n567), .Q(Address[21]) );
  FD2 Address_reg_22_ ( .D(n5505), .CP(CLOCK), .CD(n567), .Q(Address[22]) );
  FD2 Address_reg_23_ ( .D(n5506), .CP(CLOCK), .CD(n567), .Q(Address[23]) );
  FD2 Address_reg_24_ ( .D(n5507), .CP(CLOCK), .CD(n567), .Q(Address[24]) );
  FD2 Address_reg_25_ ( .D(n5508), .CP(CLOCK), .CD(n567), .Q(Address[25]) );
  FD2 Address_reg_26_ ( .D(n5509), .CP(CLOCK), .CD(n567), .Q(Address[26]) );
  FD2 Address_reg_27_ ( .D(n5510), .CP(CLOCK), .CD(n567), .Q(Address[27]) );
  FD2 Address_reg_28_ ( .D(n5511), .CP(CLOCK), .CD(n567), .Q(Address[28]) );
  FD2 Address_reg_29_ ( .D(n5512), .CP(CLOCK), .CD(n567), .Q(Address[29]) );
  FD2 ByteEnable_reg_3_ ( .D(n2910), .CP(CLOCK), .CD(n567), .QN(n4648) );
  FD2 BE_n_reg_3_ ( .D(n2909), .CP(CLOCK), .CD(n567), .Q(BE_n[3]), .QN(n5411)
         );
  FD2 ByteEnable_reg_2_ ( .D(n2908), .CP(CLOCK), .CD(n567), .QN(n4356) );
  FD2 BE_n_reg_2_ ( .D(n5523), .CP(CLOCK), .CD(n567), .Q(BE_n[2]), .QN(n5298)
         );
  FD2 ByteEnable_reg_1_ ( .D(n2907), .CP(CLOCK), .CD(n567), .QN(n4649) );
  FD2 BE_n_reg_1_ ( .D(n5522), .CP(CLOCK), .CD(n567), .Q(BE_n[1]), .QN(n5296)
         );
  FD2 ByteEnable_reg_0_ ( .D(n2906), .CP(CLOCK), .CD(n567), .QN(n4650) );
  FD2 BE_n_reg_0_ ( .D(n2905), .CP(CLOCK), .CD(n567), .Q(BE_n[0]), .QN(n5409)
         );
  ND2 U2592 ( .A(n2242), .B(n2243), .Z(n73) );
  AO7 U2593 ( .A(n2244), .B(n2245), .C(n2216), .Z(n2243) );
  IV U2594 ( .A(RESET), .Z(n567) );
  MUX21L U2595 ( .A(n5298), .B(n4356), .S(n2246), .Z(n5523) );
  MUX21L U2596 ( .A(n5296), .B(n4649), .S(n2246), .Z(n5522) );
  MUX21H U2597 ( .A(Address[0]), .B(N558), .S(n2246), .Z(n5521) );
  MUX21H U2598 ( .A(Address[3]), .B(N561), .S(n2246), .Z(n5520) );
  MUX21H U2599 ( .A(Address[2]), .B(N560), .S(n2246), .Z(n5519) );
  MUX21H U2600 ( .A(Address[5]), .B(N563), .S(n2246), .Z(n5518) );
  MUX21H U2601 ( .A(Address[4]), .B(N562), .S(n2246), .Z(n5517) );
  MUX21H U2602 ( .A(Address[7]), .B(N565), .S(n2246), .Z(n5516) );
  MUX21H U2603 ( .A(Address[6]), .B(N564), .S(n2246), .Z(n5515) );
  MUX21H U2604 ( .A(Address[9]), .B(N567), .S(n2246), .Z(n5514) );
  MUX21H U2605 ( .A(Address[8]), .B(N566), .S(n2246), .Z(n5513) );
  MUX21H U2606 ( .A(Address[29]), .B(N587), .S(n2246), .Z(n5512) );
  MUX21H U2607 ( .A(Address[28]), .B(N586), .S(n2246), .Z(n5511) );
  MUX21H U2608 ( .A(Address[27]), .B(N585), .S(n2246), .Z(n5510) );
  MUX21H U2609 ( .A(Address[26]), .B(N584), .S(n2246), .Z(n5509) );
  MUX21H U2610 ( .A(Address[25]), .B(N583), .S(n2246), .Z(n5508) );
  MUX21H U2611 ( .A(Address[24]), .B(N582), .S(n2246), .Z(n5507) );
  MUX21H U2612 ( .A(Address[23]), .B(N581), .S(n2246), .Z(n5506) );
  MUX21H U2613 ( .A(Address[22]), .B(N580), .S(n2246), .Z(n5505) );
  MUX21H U2614 ( .A(Address[21]), .B(N579), .S(n2246), .Z(n5504) );
  MUX21H U2615 ( .A(Address[20]), .B(N578), .S(n2246), .Z(n5503) );
  MUX21H U2616 ( .A(Address[19]), .B(N577), .S(n2246), .Z(n5502) );
  MUX21H U2617 ( .A(Address[18]), .B(N576), .S(n2246), .Z(n5501) );
  MUX21H U2618 ( .A(Address[17]), .B(N575), .S(n2246), .Z(n5500) );
  MUX21H U2619 ( .A(Address[16]), .B(N574), .S(n2246), .Z(n5499) );
  MUX21H U2620 ( .A(Address[15]), .B(N573), .S(n2246), .Z(n5498) );
  MUX21H U2621 ( .A(Address[14]), .B(N572), .S(n2246), .Z(n5497) );
  MUX21H U2622 ( .A(Address[13]), .B(N571), .S(n2246), .Z(n5496) );
  MUX21H U2623 ( .A(Address[12]), .B(N570), .S(n2246), .Z(n5495) );
  MUX21H U2624 ( .A(Address[11]), .B(N569), .S(n2246), .Z(n5494) );
  MUX21H U2625 ( .A(Address[10]), .B(N568), .S(n2246), .Z(n5493) );
  MUX21H U2626 ( .A(Address[1]), .B(N559), .S(n2246), .Z(n5492) );
  ND4 U2627 ( .A(n2247), .B(n2248), .C(n2249), .D(n2250), .Z(n5490) );
  NR2 U2628 ( .A(U3_U14_Z_7), .B(n2251), .Z(n2249) );
  AO2 U2629 ( .A(n2252), .B(n2253), .C(n4425), .D(n2254), .Z(n2247) );
  AO3 U2630 ( .A(n2255), .B(n2256), .C(n2257), .D(n2258), .Z(n5489) );
  MUX21L U2631 ( .A(n2259), .B(n2145), .S(n2260), .Z(n2258) );
  NR2 U2632 ( .A(n4654), .B(n2261), .Z(n2259) );
  ND2 U2633 ( .A(n2262), .B(n4468), .Z(n2257) );
  AO7 U2634 ( .A(n4458), .B(n2263), .C(n2261), .Z(n5488) );
  AO3 U2635 ( .A(n2264), .B(n2265), .C(n2266), .D(n2267), .Z(n35) );
  AO2 U2636 ( .A(n2268), .B(n2269), .C(Datai[7]), .D(n2270), .Z(n2267) );
  MUX21L U2637 ( .A(n2271), .B(n4379), .S(n2272), .Z(n2266) );
  MUX21L U2638 ( .A(n2273), .B(n4451), .S(n2274), .Z(n3287) );
  NR3 U2639 ( .A(n2275), .B(n2276), .C(n2277), .Z(n2274) );
  AO1 U2640 ( .A(n2278), .B(n2279), .C(n2280), .D(n2281), .Z(n2273) );
  IV U2641 ( .A(n2282), .Z(n2280) );
  AO3 U2642 ( .A(n2283), .B(n2284), .C(n2285), .D(n2286), .Z(n2279) );
  AO7 U2643 ( .A(n2287), .B(n4665), .C(n2288), .Z(n2285) );
  NR2 U2644 ( .A(n2289), .B(n2290), .Z(n3286) );
  NR3 U2645 ( .A(n2291), .B(n2246), .C(n2292), .Z(n2290) );
  IV U2646 ( .A(NA_n), .Z(n2291) );
  AN4 U2647 ( .A(n2293), .B(n2294), .C(n2295), .D(n2296), .Z(n2289) );
  AO3 U2648 ( .A(n2297), .B(n4451), .C(HOLD), .D(n2292), .Z(n2295) );
  OR3 U2649 ( .A(n2286), .B(n2298), .C(n2299), .Z(n2293) );
  AO3 U2650 ( .A(n4451), .B(n2300), .C(n2296), .D(n2301), .Z(n3285) );
  AO1 U2651 ( .A(n2297), .B(n2302), .C(n2303), .D(n2304), .Z(n2301) );
  AO6 U2652 ( .A(n2298), .B(n2286), .C(n2305), .Z(n2304) );
  IV U2653 ( .A(n2306), .Z(n2305) );
  NR2 U2654 ( .A(n2217), .B(HOLD), .Z(n2298) );
  IV U2655 ( .A(n2307), .Z(n2303) );
  AO6 U2656 ( .A(n2308), .B(READY_n), .C(n2309), .Z(n2296) );
  ND4 U2657 ( .A(n2307), .B(n2299), .C(n2310), .D(n2311), .Z(n3284) );
  AO2 U2658 ( .A(n4451), .B(n2292), .C(n2297), .D(HOLD), .Z(n2311) );
  IV U2659 ( .A(n2312), .Z(n2297) );
  ND2 U2660 ( .A(n2312), .B(n2300), .Z(n2292) );
  ND3 U2661 ( .A(n4667), .B(n4651), .C(n4666), .Z(n2300) );
  ND2 U2662 ( .A(n4666), .B(n2184), .Z(n2312) );
  AO7 U2663 ( .A(READY_n), .B(n2313), .C(n2306), .Z(n2299) );
  ND2 U2664 ( .A(n2284), .B(n2314), .Z(n2307) );
  OR3 U2665 ( .A(n2315), .B(NA_n), .C(n2313), .Z(n2314) );
  IV U2666 ( .A(n2302), .Z(n2313) );
  NR2 U2667 ( .A(HOLD), .B(n4451), .Z(n2302) );
  AO7 U2668 ( .A(n5397), .B(n2246), .C(n2316), .Z(n3283) );
  AO7 U2669 ( .A(n4665), .B(n2317), .C(n2318), .Z(n3282) );
  AO4 U2670 ( .A(n4655), .B(n2317), .C(BS16_n), .D(n2319), .Z(n3281) );
  AO7 U2671 ( .A(n4656), .B(n2317), .C(n2318), .Z(n3280) );
  AO6 U2672 ( .A(n2320), .B(BS16_n), .C(n2321), .Z(n2318) );
  IV U2673 ( .A(n2316), .Z(n2317) );
  NR2 U2674 ( .A(n2320), .B(n2321), .Z(n2316) );
  IV U2675 ( .A(n2319), .Z(n2320) );
  NR2 U2676 ( .A(n2309), .B(n2306), .Z(n2319) );
  AN3 U2677 ( .A(n4651), .B(n2150), .C(n4666), .Z(n2306) );
  AO3 U2678 ( .A(n4647), .B(n2322), .C(n2323), .D(n2324), .Z(n3279) );
  AO6 U2679 ( .A(n203), .B(n2325), .C(n2326), .Z(n2324) );
  AO4 U2680 ( .A(n2327), .B(n2328), .C(n4646), .D(n2329), .Z(n2326) );
  AO2 U2681 ( .A(n429), .B(n2330), .C(rEIP[31]), .D(n2331), .Z(n2323) );
  AO3 U2682 ( .A(n2328), .B(n2332), .C(n2333), .D(n2334), .Z(n3278) );
  AO2 U2683 ( .A(n429), .B(n2276), .C(n2335), .D(rEIP[31]), .Z(n2334) );
  OR2 U2684 ( .A(n2336), .B(n4647), .Z(n2333) );
  IV U2685 ( .A(n286), .Z(n2328) );
  AO3 U2686 ( .A(n2337), .B(n2338), .C(n2339), .D(n2340), .Z(n3277) );
  AO2 U2687 ( .A(n2341), .B(n4657), .C(n2335), .D(rEIP[31]), .Z(n2340) );
  ND2 U2688 ( .A(n2342), .B(n286), .Z(n2339) );
  AO7 U2689 ( .A(n4467), .B(n2343), .C(n2344), .Z(n3276) );
  EO1 U2690 ( .A(n2262), .B(n2345), .C(n2256), .D(n2346), .Z(n2344) );
  AO7 U2691 ( .A(n2347), .B(n2348), .C(n2349), .Z(n2345) );
  IV U2692 ( .A(n2350), .Z(n2343) );
  MUX21L U2693 ( .A(n4658), .B(n2351), .S(n2263), .Z(n3275) );
  AO1 U2694 ( .A(n2352), .B(n2353), .C(n2354), .D(n2355), .Z(n2351) );
  ND2 U2695 ( .A(n2356), .B(n2357), .Z(n2354) );
  AO7 U2696 ( .A(n2281), .B(n2358), .C(READY_n), .Z(n2356) );
  ND4 U2697 ( .A(n2359), .B(n2360), .C(n2357), .D(n2361), .Z(n3274) );
  AO1 U2698 ( .A(n2362), .B(n2170), .C(n2363), .D(n2364), .Z(n2361) );
  NR2 U2699 ( .A(READY_n), .B(n2365), .Z(n2363) );
  MUX21L U2700 ( .A(n4668), .B(n2366), .S(n2263), .Z(n3273) );
  IV U2701 ( .A(n2362), .Z(n2263) );
  NR3 U2702 ( .A(n2277), .B(n2355), .C(n2367), .Z(n2362) );
  AO3 U2703 ( .A(n2359), .B(n2368), .C(n2261), .D(n2242), .Z(n2367) );
  AO3 U2704 ( .A(n2369), .B(n2359), .C(n2322), .D(n2370), .Z(n2355) );
  AO1 U2705 ( .A(n2371), .B(n2372), .C(n2373), .D(n2374), .Z(n2369) );
  AO4 U2706 ( .A(n2346), .B(n2375), .C(n2376), .D(n2171), .Z(n2374) );
  AN2 U2707 ( .A(n2375), .B(n2346), .Z(n2376) );
  AO7 U2708 ( .A(n4456), .B(n2377), .C(n2378), .Z(n2375) );
  AO4 U2709 ( .A(n2379), .B(n2380), .C(n2147), .D(n2381), .Z(n2378) );
  AO1 U2710 ( .A(n4455), .B(n2382), .C(n2383), .D(n4454), .Z(n2380) );
  IV U2711 ( .A(n2255), .Z(n2383) );
  EN U2712 ( .A(n4468), .B(n2384), .Z(n2255) );
  NR2 U2713 ( .A(n4455), .B(n2382), .Z(n2379) );
  AO3 U2714 ( .A(n2385), .B(n2386), .C(n2387), .D(n2353), .Z(n2373) );
  AN2 U2715 ( .A(n4357), .B(n4355), .Z(n2385) );
  AO7 U2716 ( .A(READY_n), .B(n2357), .C(n2365), .Z(n2277) );
  NR3 U2717 ( .A(n2388), .B(n2278), .C(n2389), .Z(n2366) );
  MUX21L U2718 ( .A(n2242), .B(n2365), .S(READY_n), .Z(n2388) );
  IV U2719 ( .A(n2281), .Z(n2365) );
  AN3 U2720 ( .A(n4450), .B(n2151), .C(n2390), .Z(n2281) );
  MUX21L U2721 ( .A(n2215), .B(n2391), .S(n2275), .Z(n3272) );
  NR2 U2722 ( .A(n2392), .B(n2393), .Z(n2391) );
  MUX21L U2723 ( .A(n5430), .B(n4354), .S(n2246), .Z(n3271) );
  MUX21L U2724 ( .A(n4462), .B(n2394), .S(n2275), .Z(n3270) );
  AO7 U2725 ( .A(n2244), .B(n2245), .C(n2282), .Z(n2275) );
  NR2 U2726 ( .A(n2288), .B(n2393), .Z(n2394) );
  ND2 U2727 ( .A(n2282), .B(n2395), .Z(n2393) );
  NR2 U2728 ( .A(n2335), .B(n2358), .Z(n2282) );
  IV U2729 ( .A(n2242), .Z(n2358) );
  OR3 U2730 ( .A(n4658), .B(n2396), .C(n2170), .Z(n2242) );
  MUX21L U2731 ( .A(n5429), .B(n4462), .S(n2246), .Z(n3269) );
  AO3 U2732 ( .A(n4460), .B(n2322), .C(n2397), .D(n2398), .Z(n3268) );
  IV U2733 ( .A(n2399), .Z(n2398) );
  AO3 U2734 ( .A(n2329), .B(n4463), .C(n2400), .D(n2401), .Z(n2399) );
  ND2 U2735 ( .A(n2402), .B(N2787), .Z(n2401) );
  AO2 U2736 ( .A(n2325), .B(n234), .C(n2403), .D(n317), .Z(n2400) );
  AO2 U2737 ( .A(n460), .B(n2330), .C(rEIP[0]), .D(n2331), .Z(n2397) );
  AO3 U2738 ( .A(n4459), .B(n2322), .C(n2404), .D(n2405), .Z(n3267) );
  IV U2739 ( .A(n2406), .Z(n2405) );
  AO3 U2740 ( .A(n2329), .B(n4452), .C(n2407), .D(n2408), .Z(n2406) );
  ND2 U2741 ( .A(n2402), .B(N2788), .Z(n2408) );
  AO2 U2742 ( .A(n2325), .B(n233), .C(n2403), .D(n316), .Z(n2407) );
  AO2 U2743 ( .A(n459), .B(n2330), .C(rEIP[1]), .D(n2331), .Z(n2404) );
  AO3 U2744 ( .A(n4472), .B(n2322), .C(n2409), .D(n2410), .Z(n3266) );
  IV U2745 ( .A(n2411), .Z(n2410) );
  AO3 U2746 ( .A(n2329), .B(n4471), .C(n2412), .D(n2413), .Z(n2411) );
  ND2 U2747 ( .A(n2402), .B(N2789), .Z(n2413) );
  AO2 U2748 ( .A(n2325), .B(n232), .C(n2403), .D(n315), .Z(n2412) );
  AO2 U2749 ( .A(n458), .B(n2330), .C(rEIP[2]), .D(n2331), .Z(n2409) );
  AO3 U2750 ( .A(n4477), .B(n2322), .C(n2414), .D(n2415), .Z(n3265) );
  IV U2751 ( .A(n2416), .Z(n2415) );
  AO3 U2752 ( .A(n2329), .B(n4476), .C(n2417), .D(n2418), .Z(n2416) );
  ND2 U2753 ( .A(n2402), .B(N2790), .Z(n2418) );
  AO2 U2754 ( .A(n2325), .B(n231), .C(n2403), .D(n314), .Z(n2417) );
  AO2 U2755 ( .A(n457), .B(n2330), .C(rEIP[3]), .D(n2331), .Z(n2414) );
  ND4 U2756 ( .A(n2419), .B(n2420), .C(n2421), .D(n2422), .Z(n3264) );
  AO6 U2757 ( .A(N2791), .B(n2402), .C(n2335), .Z(n2422) );
  EO1 U2758 ( .A(n313), .B(n2403), .C(n2329), .D(n4481), .Z(n2421) );
  AO2 U2759 ( .A(n230), .B(n2325), .C(n456), .D(n2330), .Z(n2420) );
  AO2 U2760 ( .A(rEIP[4]), .B(n2331), .C(n2423), .D(n2185), .Z(n2419) );
  ND4 U2761 ( .A(n2424), .B(n2425), .C(n2426), .D(n2427), .Z(n3263) );
  AO6 U2762 ( .A(N2792), .B(n2402), .C(n2335), .Z(n2427) );
  NR2 U2763 ( .A(n2428), .B(n2429), .Z(n2402) );
  EO1 U2764 ( .A(n312), .B(n2403), .C(n2329), .D(n4486), .Z(n2426) );
  IV U2765 ( .A(n2327), .Z(n2403) );
  AO2 U2766 ( .A(n229), .B(n2325), .C(n455), .D(n2330), .Z(n2425) );
  AO2 U2767 ( .A(rEIP[5]), .B(n2331), .C(n2423), .D(n2186), .Z(n2424) );
  AO3 U2768 ( .A(n4492), .B(n2322), .C(n2430), .D(n2431), .Z(n3262) );
  AO1 U2769 ( .A(n2432), .B(n2218), .C(n2433), .D(n2335), .Z(n2431) );
  AO4 U2770 ( .A(n2434), .B(n2435), .C(n2327), .D(n2436), .Z(n2433) );
  AO2 U2771 ( .A(n454), .B(n2330), .C(rEIP[6]), .D(n2331), .Z(n2430) );
  AO3 U2772 ( .A(n4497), .B(n2322), .C(n2437), .D(n2438), .Z(n3261) );
  AO1 U2773 ( .A(n2432), .B(n2219), .C(n2439), .D(n2335), .Z(n2438) );
  AO4 U2774 ( .A(n2434), .B(n2440), .C(n2327), .D(n2441), .Z(n2439) );
  AO2 U2775 ( .A(n453), .B(n2330), .C(rEIP[7]), .D(n2331), .Z(n2437) );
  AO3 U2776 ( .A(n4502), .B(n2322), .C(n2442), .D(n2443), .Z(n3260) );
  AO1 U2777 ( .A(n2432), .B(n2220), .C(n2444), .D(n2335), .Z(n2443) );
  AO4 U2778 ( .A(n2434), .B(n2445), .C(n2327), .D(n2446), .Z(n2444) );
  AO2 U2779 ( .A(n452), .B(n2330), .C(rEIP[8]), .D(n2331), .Z(n2442) );
  AO3 U2780 ( .A(n4506), .B(n2322), .C(n2447), .D(n2448), .Z(n3259) );
  AO1 U2781 ( .A(n2432), .B(n2221), .C(n2449), .D(n2335), .Z(n2448) );
  AO4 U2782 ( .A(n2434), .B(n2450), .C(n2327), .D(n2451), .Z(n2449) );
  AO2 U2783 ( .A(n451), .B(n2330), .C(rEIP[9]), .D(n2331), .Z(n2447) );
  AO3 U2784 ( .A(n4510), .B(n2322), .C(n2452), .D(n2453), .Z(n3258) );
  AO1 U2785 ( .A(n2432), .B(n2222), .C(n2454), .D(n2335), .Z(n2453) );
  AO4 U2786 ( .A(n2434), .B(n2455), .C(n2327), .D(n2456), .Z(n2454) );
  AO2 U2787 ( .A(n450), .B(n2330), .C(rEIP[10]), .D(n2331), .Z(n2452) );
  AO3 U2788 ( .A(n4514), .B(n2322), .C(n2457), .D(n2458), .Z(n3257) );
  AO1 U2789 ( .A(n2432), .B(n2223), .C(n2459), .D(n2335), .Z(n2458) );
  AO4 U2790 ( .A(n2434), .B(n2460), .C(n2327), .D(n2461), .Z(n2459) );
  AO2 U2791 ( .A(n449), .B(n2330), .C(rEIP[11]), .D(n2331), .Z(n2457) );
  AO3 U2792 ( .A(n4518), .B(n2322), .C(n2462), .D(n2463), .Z(n3256) );
  AO1 U2793 ( .A(n2432), .B(n2224), .C(n2464), .D(n2335), .Z(n2463) );
  AO4 U2794 ( .A(n2434), .B(n2465), .C(n2327), .D(n2466), .Z(n2464) );
  AO2 U2795 ( .A(n448), .B(n2330), .C(rEIP[12]), .D(n2331), .Z(n2462) );
  AO3 U2796 ( .A(n4522), .B(n2322), .C(n2467), .D(n2468), .Z(n3255) );
  AO1 U2797 ( .A(n2432), .B(n2225), .C(n2469), .D(n2335), .Z(n2468) );
  AO4 U2798 ( .A(n2434), .B(n2470), .C(n2327), .D(n2471), .Z(n2469) );
  AO2 U2799 ( .A(n447), .B(n2330), .C(rEIP[13]), .D(n2331), .Z(n2467) );
  AO3 U2800 ( .A(n4526), .B(n2322), .C(n2472), .D(n2473), .Z(n3254) );
  AO1 U2801 ( .A(n2432), .B(n2226), .C(n2474), .D(n2335), .Z(n2473) );
  AO4 U2802 ( .A(n2434), .B(n2475), .C(n2327), .D(n2476), .Z(n2474) );
  AO2 U2803 ( .A(n446), .B(n2330), .C(rEIP[14]), .D(n2331), .Z(n2472) );
  AO3 U2804 ( .A(n4530), .B(n2322), .C(n2477), .D(n2478), .Z(n3253) );
  AO1 U2805 ( .A(n2432), .B(n2227), .C(n2479), .D(n2335), .Z(n2478) );
  AO4 U2806 ( .A(n2434), .B(n2480), .C(n2327), .D(n2481), .Z(n2479) );
  AO2 U2807 ( .A(n445), .B(n2330), .C(rEIP[15]), .D(n2331), .Z(n2477) );
  AO3 U2808 ( .A(n4535), .B(n2322), .C(n2482), .D(n2483), .Z(n3252) );
  AO1 U2809 ( .A(n2432), .B(n2190), .C(n2484), .D(n2335), .Z(n2483) );
  AO4 U2810 ( .A(n2434), .B(n2485), .C(n2327), .D(n2486), .Z(n2484) );
  AO2 U2811 ( .A(n444), .B(n2330), .C(rEIP[16]), .D(n2331), .Z(n2482) );
  AO3 U2812 ( .A(n4539), .B(n2322), .C(n2487), .D(n2488), .Z(n3251) );
  AO1 U2813 ( .A(n2432), .B(n2189), .C(n2489), .D(n2335), .Z(n2488) );
  AO4 U2814 ( .A(n2434), .B(n2490), .C(n2327), .D(n2491), .Z(n2489) );
  AO2 U2815 ( .A(n443), .B(n2330), .C(rEIP[17]), .D(n2331), .Z(n2487) );
  AO3 U2816 ( .A(n4543), .B(n2322), .C(n2492), .D(n2493), .Z(n3250) );
  AO1 U2817 ( .A(n2432), .B(n2188), .C(n2494), .D(n2335), .Z(n2493) );
  AO4 U2818 ( .A(n2434), .B(n2495), .C(n2327), .D(n2496), .Z(n2494) );
  AO2 U2819 ( .A(n442), .B(n2330), .C(rEIP[18]), .D(n2331), .Z(n2492) );
  AO3 U2820 ( .A(n4547), .B(n2322), .C(n2497), .D(n2498), .Z(n3249) );
  AO1 U2821 ( .A(n2432), .B(n2187), .C(n2499), .D(n2335), .Z(n2498) );
  AO4 U2822 ( .A(n2434), .B(n2500), .C(n2327), .D(n2501), .Z(n2499) );
  IV U2823 ( .A(n2329), .Z(n2432) );
  AO2 U2824 ( .A(n441), .B(n2330), .C(rEIP[19]), .D(n2331), .Z(n2497) );
  AO3 U2825 ( .A(n4551), .B(n2322), .C(n2502), .D(n2503), .Z(n3248) );
  AO6 U2826 ( .A(n214), .B(n2325), .C(n2504), .Z(n2503) );
  AO4 U2827 ( .A(n2327), .B(n2505), .C(n4550), .D(n2329), .Z(n2504) );
  AO2 U2828 ( .A(n440), .B(n2330), .C(rEIP[20]), .D(n2331), .Z(n2502) );
  AO3 U2829 ( .A(n4555), .B(n2322), .C(n2506), .D(n2507), .Z(n3247) );
  AO6 U2830 ( .A(n213), .B(n2325), .C(n2508), .Z(n2507) );
  AO4 U2831 ( .A(n2327), .B(n2509), .C(n4554), .D(n2329), .Z(n2508) );
  AO2 U2832 ( .A(n439), .B(n2330), .C(rEIP[21]), .D(n2331), .Z(n2506) );
  AO3 U2833 ( .A(n4559), .B(n2322), .C(n2510), .D(n2511), .Z(n3246) );
  AO6 U2834 ( .A(n212), .B(n2325), .C(n2512), .Z(n2511) );
  AO4 U2835 ( .A(n2327), .B(n2513), .C(n4558), .D(n2329), .Z(n2512) );
  AO2 U2836 ( .A(n438), .B(n2330), .C(rEIP[22]), .D(n2331), .Z(n2510) );
  AO3 U2837 ( .A(n4563), .B(n2322), .C(n2514), .D(n2515), .Z(n3245) );
  AO6 U2838 ( .A(n211), .B(n2325), .C(n2516), .Z(n2515) );
  AO4 U2839 ( .A(n2327), .B(n2517), .C(n4562), .D(n2329), .Z(n2516) );
  AO2 U2840 ( .A(n437), .B(n2330), .C(rEIP[23]), .D(n2331), .Z(n2514) );
  AO3 U2841 ( .A(n4567), .B(n2322), .C(n2518), .D(n2519), .Z(n3244) );
  AO6 U2842 ( .A(n210), .B(n2325), .C(n2520), .Z(n2519) );
  AO4 U2843 ( .A(n2327), .B(n2521), .C(n4566), .D(n2329), .Z(n2520) );
  AO2 U2844 ( .A(n436), .B(n2330), .C(rEIP[24]), .D(n2331), .Z(n2518) );
  AO3 U2845 ( .A(n4571), .B(n2322), .C(n2522), .D(n2523), .Z(n3243) );
  AO6 U2846 ( .A(n209), .B(n2325), .C(n2524), .Z(n2523) );
  AO4 U2847 ( .A(n2327), .B(n2525), .C(n4570), .D(n2329), .Z(n2524) );
  AO2 U2848 ( .A(n435), .B(n2330), .C(rEIP[25]), .D(n2331), .Z(n2522) );
  AO3 U2849 ( .A(n4575), .B(n2322), .C(n2526), .D(n2527), .Z(n3242) );
  AO6 U2850 ( .A(n208), .B(n2325), .C(n2528), .Z(n2527) );
  AO4 U2851 ( .A(n2327), .B(n2529), .C(n4574), .D(n2329), .Z(n2528) );
  AO2 U2852 ( .A(n434), .B(n2330), .C(rEIP[26]), .D(n2331), .Z(n2526) );
  AO3 U2853 ( .A(n4579), .B(n2322), .C(n2530), .D(n2531), .Z(n3241) );
  AO6 U2854 ( .A(n207), .B(n2325), .C(n2532), .Z(n2531) );
  AO4 U2855 ( .A(n2327), .B(n2533), .C(n4578), .D(n2329), .Z(n2532) );
  AO2 U2856 ( .A(n433), .B(n2330), .C(rEIP[27]), .D(n2331), .Z(n2530) );
  AO3 U2857 ( .A(n4583), .B(n2322), .C(n2534), .D(n2535), .Z(n3240) );
  AO6 U2858 ( .A(n206), .B(n2325), .C(n2536), .Z(n2535) );
  AO4 U2859 ( .A(n2327), .B(n2537), .C(n4582), .D(n2329), .Z(n2536) );
  AO2 U2860 ( .A(n432), .B(n2330), .C(rEIP[28]), .D(n2331), .Z(n2534) );
  AO3 U2861 ( .A(n4587), .B(n2322), .C(n2538), .D(n2539), .Z(n3239) );
  AO6 U2862 ( .A(n205), .B(n2325), .C(n2540), .Z(n2539) );
  AO4 U2863 ( .A(n2327), .B(n2541), .C(n4586), .D(n2329), .Z(n2540) );
  AO2 U2864 ( .A(n431), .B(n2330), .C(rEIP[29]), .D(n2331), .Z(n2538) );
  AO3 U2865 ( .A(n4644), .B(n2322), .C(n2542), .D(n2543), .Z(n3238) );
  AO6 U2866 ( .A(n204), .B(n2325), .C(n2544), .Z(n2543) );
  AO4 U2867 ( .A(n2327), .B(n2545), .C(n4643), .D(n2329), .Z(n2544) );
  ND2 U2868 ( .A(n2546), .B(n2547), .Z(n2329) );
  AO4 U2869 ( .A(n2548), .B(n2549), .C(n2550), .D(n2551), .Z(n2547) );
  ND2 U2870 ( .A(n2552), .B(n2553), .Z(n2551) );
  ND3 U2871 ( .A(n2288), .B(n2548), .C(n2546), .Z(n2327) );
  IV U2872 ( .A(n2434), .Z(n2325) );
  ND2 U2873 ( .A(n2550), .B(n2554), .Z(n2434) );
  AO7 U2874 ( .A(n2555), .B(n2428), .C(n2556), .Z(n2554) );
  AO2 U2875 ( .A(n430), .B(n2330), .C(rEIP[30]), .D(n2331), .Z(n2542) );
  AO4 U2876 ( .A(n2550), .B(n2557), .C(n2428), .D(n2558), .Z(n2330) );
  ND2 U2877 ( .A(n2552), .B(n2555), .Z(n2558) );
  IV U2878 ( .A(n2553), .Z(n2555) );
  IV U2879 ( .A(n2546), .Z(n2428) );
  NR2 U2880 ( .A(n2359), .B(n2331), .Z(n2546) );
  OR2 U2881 ( .A(n2556), .B(n2331), .Z(n2557) );
  NR4 U2882 ( .A(n2559), .B(n2389), .C(n2423), .D(n2335), .Z(n2331) );
  IV U2883 ( .A(n2322), .Z(n2423) );
  NR2 U2884 ( .A(n2245), .B(n2244), .Z(n2559) );
  ND4 U2885 ( .A(n4450), .B(n4668), .C(n2151), .D(n2183), .Z(n2322) );
  ND2 U2886 ( .A(n2560), .B(n2310), .Z(n3236) );
  IV U2887 ( .A(n2321), .Z(n2310) );
  NR3 U2888 ( .A(n2184), .B(n4666), .C(n2150), .Z(n2321) );
  MUX21L U2889 ( .A(D_C_n), .B(n4652), .S(n2246), .Z(n2560) );
  AO3 U2890 ( .A(n2561), .B(n2562), .C(n2563), .D(n2564), .Z(n3234) );
  AO2 U2891 ( .A(n2565), .B(n2382), .C(n2260), .D(n2167), .Z(n2564) );
  IV U2892 ( .A(n2566), .Z(n2260) );
  EO U2893 ( .A(n2567), .B(n2568), .Z(n2382) );
  ND2 U2894 ( .A(n2569), .B(n2570), .Z(n2568) );
  MUX21L U2895 ( .A(n2167), .B(n2571), .S(n2572), .Z(n2569) );
  IV U2896 ( .A(n2256), .Z(n2565) );
  AO7 U2897 ( .A(n2573), .B(n2571), .C(n2262), .Z(n2563) );
  AO3 U2898 ( .A(n2256), .B(n2381), .C(n2574), .D(n2575), .Z(n3233) );
  MUX21L U2899 ( .A(n2350), .B(n2576), .S(n4653), .Z(n2575) );
  NR2 U2900 ( .A(n2348), .B(n2577), .Z(n2576) );
  AO7 U2901 ( .A(n2578), .B(n2577), .C(n2566), .Z(n2350) );
  ND2 U2902 ( .A(n2561), .B(n2579), .Z(n2574) );
  IV U2903 ( .A(n2562), .Z(n2579) );
  ND3 U2904 ( .A(n2352), .B(n2566), .C(n4654), .Z(n2562) );
  EO U2905 ( .A(n4453), .B(n2550), .Z(n2561) );
  ND2 U2906 ( .A(n2278), .B(n2566), .Z(n2256) );
  OR3 U2907 ( .A(n2580), .B(n2262), .C(n2581), .Z(n2566) );
  ND2 U2908 ( .A(n2582), .B(n2583), .Z(n3231) );
  ND3 U2909 ( .A(n2584), .B(n2353), .C(n2352), .Z(n2583) );
  MUX21L U2910 ( .A(n2585), .B(n2262), .S(n4454), .Z(n2582) );
  AO3 U2911 ( .A(n2586), .B(n2262), .C(n2584), .D(n2556), .Z(n2585) );
  AO7 U2912 ( .A(n2586), .B(n2587), .C(n2588), .Z(n3230) );
  MUX21L U2913 ( .A(n2589), .B(n2389), .S(n4455), .Z(n2588) );
  ND2 U2914 ( .A(n2590), .B(n2584), .Z(n2589) );
  EN U2915 ( .A(n2591), .B(n2592), .Z(n2587) );
  ND2 U2916 ( .A(n2593), .B(n2594), .Z(n3229) );
  MUX21L U2917 ( .A(n2595), .B(n2596), .S(n2597), .Z(n2594) );
  EO U2918 ( .A(n4456), .B(n4665), .Z(n2597) );
  AO7 U2919 ( .A(n2146), .B(n2556), .C(n2590), .Z(n2596) );
  NR2 U2920 ( .A(n4455), .B(n2598), .Z(n2595) );
  MUX21L U2921 ( .A(n2599), .B(n2600), .S(n4456), .Z(n2593) );
  AO4 U2922 ( .A(n2601), .B(n2602), .C(n4457), .D(n2603), .Z(n3228) );
  AO1 U2923 ( .A(n2389), .B(n4455), .C(n2599), .D(n2604), .Z(n2603) );
  AO6 U2924 ( .A(n2586), .B(n2556), .C(n2147), .Z(n2604) );
  AO7 U2925 ( .A(n2586), .B(n2600), .C(n2584), .Z(n2599) );
  AO3 U2926 ( .A(n2261), .B(n2353), .C(n2605), .D(n2606), .Z(n2584) );
  IV U2927 ( .A(n2581), .Z(n2605) );
  ND2 U2928 ( .A(n2607), .B(n2608), .Z(n2353) );
  AO7 U2929 ( .A(n2359), .B(n2381), .C(n2609), .Z(n2608) );
  ND4 U2930 ( .A(n4357), .B(n2352), .C(n2610), .D(n2148), .Z(n2609) );
  IV U2931 ( .A(n2377), .Z(n2381) );
  EO U2932 ( .A(n2611), .B(n2612), .Z(n2377) );
  EO U2933 ( .A(n4653), .B(n2613), .Z(n2612) );
  AO4 U2934 ( .A(n4467), .B(n2261), .C(n2346), .D(n2359), .Z(n2607) );
  EO U2935 ( .A(n4467), .B(n2614), .Z(n2346) );
  AO5 U2936 ( .A(n2615), .B(n4653), .C(n2611), .Z(n2614) );
  AO2 U2937 ( .A(n2167), .B(n2567), .C(n2578), .D(n2572), .Z(n2611) );
  IV U2938 ( .A(n2384), .Z(n2572) );
  ND2 U2939 ( .A(n2244), .B(n2250), .Z(n2384) );
  ND3 U2940 ( .A(n2616), .B(n2250), .C(n2248), .Z(n2567) );
  NR2 U2941 ( .A(n2262), .B(n2617), .Z(n2586) );
  AO1 U2942 ( .A(n2618), .B(n2146), .C(n2600), .D(n2364), .Z(n2601) );
  AO4 U2943 ( .A(n4455), .B(n2360), .C(n2592), .D(n2591), .Z(n2600) );
  ND2 U2944 ( .A(n2262), .B(n2169), .Z(n2591) );
  EO U2945 ( .A(n2146), .B(n2360), .Z(n2592) );
  AO3 U2946 ( .A(n2619), .B(n2620), .C(n2621), .D(n2622), .Z(n3227) );
  AO2 U2947 ( .A(n2623), .B(n445), .C(n4531), .D(n2624), .Z(n2622) );
  ND2 U2948 ( .A(N2594), .B(n2625), .Z(n2621) );
  AO7 U2949 ( .A(n4466), .B(n2626), .C(n2627), .Z(n3226) );
  AO2 U2950 ( .A(Datai[0]), .B(n2628), .C(n4465), .D(n2629), .Z(n2627) );
  AO7 U2951 ( .A(n4470), .B(n2626), .C(n2630), .Z(n3225) );
  AO2 U2952 ( .A(Datai[1]), .B(n2628), .C(n4469), .D(n2629), .Z(n2630) );
  AO7 U2953 ( .A(n4475), .B(n2626), .C(n2631), .Z(n3224) );
  AO2 U2954 ( .A(Datai[2]), .B(n2628), .C(n4474), .D(n2629), .Z(n2631) );
  AO7 U2955 ( .A(n4480), .B(n2626), .C(n2632), .Z(n3223) );
  AO2 U2956 ( .A(Datai[3]), .B(n2628), .C(n4479), .D(n2629), .Z(n2632) );
  AO7 U2957 ( .A(n4485), .B(n2626), .C(n2633), .Z(n3222) );
  AO2 U2958 ( .A(Datai[4]), .B(n2628), .C(n4484), .D(n2629), .Z(n2633) );
  AO7 U2959 ( .A(n4490), .B(n2626), .C(n2634), .Z(n3221) );
  AO2 U2960 ( .A(Datai[5]), .B(n2628), .C(n4489), .D(n2629), .Z(n2634) );
  AO7 U2961 ( .A(n4495), .B(n2626), .C(n2635), .Z(n3220) );
  AO2 U2962 ( .A(Datai[6]), .B(n2628), .C(n4494), .D(n2629), .Z(n2635) );
  AO7 U2963 ( .A(n4500), .B(n2626), .C(n2636), .Z(n3219) );
  AO2 U2964 ( .A(n2628), .B(Datai[7]), .C(n4499), .D(n2629), .Z(n2636) );
  AO7 U2965 ( .A(n4504), .B(n2626), .C(n2637), .Z(n3218) );
  AO2 U2966 ( .A(Datai[8]), .B(n2628), .C(n4503), .D(n2629), .Z(n2637) );
  AO7 U2967 ( .A(n4508), .B(n2626), .C(n2638), .Z(n3217) );
  AO2 U2968 ( .A(Datai[9]), .B(n2628), .C(n4507), .D(n2629), .Z(n2638) );
  AO7 U2969 ( .A(n4512), .B(n2626), .C(n2639), .Z(n3216) );
  AO2 U2970 ( .A(Datai[10]), .B(n2628), .C(n4511), .D(n2629), .Z(n2639) );
  AO7 U2971 ( .A(n4516), .B(n2626), .C(n2640), .Z(n3215) );
  AO2 U2972 ( .A(Datai[11]), .B(n2628), .C(n4515), .D(n2629), .Z(n2640) );
  AO7 U2973 ( .A(n4520), .B(n2626), .C(n2641), .Z(n3214) );
  AO2 U2974 ( .A(Datai[12]), .B(n2628), .C(n4519), .D(n2629), .Z(n2641) );
  AO7 U2975 ( .A(n4524), .B(n2626), .C(n2642), .Z(n3213) );
  AO2 U2976 ( .A(Datai[13]), .B(n2628), .C(n4523), .D(n2629), .Z(n2642) );
  AO7 U2977 ( .A(n4528), .B(n2626), .C(n2643), .Z(n3212) );
  AO2 U2978 ( .A(Datai[14]), .B(n2628), .C(n4527), .D(n2629), .Z(n2643) );
  AO7 U2979 ( .A(n4532), .B(n2626), .C(n2644), .Z(n3211) );
  AO2 U2980 ( .A(n2628), .B(Datai[15]), .C(n2629), .D(n4531), .Z(n2644) );
  AO3 U2981 ( .A(n2619), .B(n2645), .C(n2646), .D(n2647), .Z(n3210) );
  AO2 U2982 ( .A(n2623), .B(n460), .C(n4465), .D(n2624), .Z(n2647) );
  ND2 U2983 ( .A(N2579), .B(n2625), .Z(n2646) );
  AO3 U2984 ( .A(n2619), .B(n2648), .C(n2649), .D(n2650), .Z(n3209) );
  AO2 U2985 ( .A(n2623), .B(n459), .C(n4469), .D(n2624), .Z(n2650) );
  ND2 U2986 ( .A(N2580), .B(n2625), .Z(n2649) );
  AO3 U2987 ( .A(n2619), .B(n2651), .C(n2652), .D(n2653), .Z(n3208) );
  AO2 U2988 ( .A(n2623), .B(n458), .C(n4474), .D(n2624), .Z(n2653) );
  ND2 U2989 ( .A(N2581), .B(n2625), .Z(n2652) );
  AO3 U2990 ( .A(n2619), .B(n2654), .C(n2655), .D(n2656), .Z(n3207) );
  AO2 U2991 ( .A(n2623), .B(n457), .C(n4479), .D(n2624), .Z(n2656) );
  ND2 U2992 ( .A(N2582), .B(n2625), .Z(n2655) );
  AO3 U2993 ( .A(n2619), .B(n2657), .C(n2658), .D(n2659), .Z(n3206) );
  AO2 U2994 ( .A(n2623), .B(n456), .C(n4484), .D(n2624), .Z(n2659) );
  ND2 U2995 ( .A(N2583), .B(n2625), .Z(n2658) );
  AO3 U2996 ( .A(n2619), .B(n2660), .C(n2661), .D(n2662), .Z(n3205) );
  AO2 U2997 ( .A(n2623), .B(n455), .C(n4489), .D(n2624), .Z(n2662) );
  ND2 U2998 ( .A(N2584), .B(n2625), .Z(n2661) );
  AO3 U2999 ( .A(n2619), .B(n2663), .C(n2664), .D(n2665), .Z(n3204) );
  AO2 U3000 ( .A(n2623), .B(n454), .C(n4494), .D(n2624), .Z(n2665) );
  ND2 U3001 ( .A(N2585), .B(n2625), .Z(n2664) );
  AO3 U3002 ( .A(n2666), .B(n2619), .C(n2667), .D(n2668), .Z(n3203) );
  AO2 U3003 ( .A(n2623), .B(n453), .C(n4499), .D(n2624), .Z(n2668) );
  ND2 U3004 ( .A(N2586), .B(n2625), .Z(n2667) );
  AO3 U3005 ( .A(n2619), .B(n2669), .C(n2670), .D(n2671), .Z(n3202) );
  AO2 U3006 ( .A(n2623), .B(n452), .C(n4503), .D(n2624), .Z(n2671) );
  ND2 U3007 ( .A(N2587), .B(n2625), .Z(n2670) );
  AO3 U3008 ( .A(n2619), .B(n2672), .C(n2673), .D(n2674), .Z(n3201) );
  AO2 U3009 ( .A(n2623), .B(n451), .C(n4507), .D(n2624), .Z(n2674) );
  ND2 U3010 ( .A(N2588), .B(n2625), .Z(n2673) );
  AO3 U3011 ( .A(n2619), .B(n2675), .C(n2676), .D(n2677), .Z(n3200) );
  AO2 U3012 ( .A(n2623), .B(n450), .C(n4511), .D(n2624), .Z(n2677) );
  ND2 U3013 ( .A(N2589), .B(n2625), .Z(n2676) );
  AO3 U3014 ( .A(n2619), .B(n2678), .C(n2679), .D(n2680), .Z(n3199) );
  AO2 U3015 ( .A(n2623), .B(n449), .C(n4515), .D(n2624), .Z(n2680) );
  ND2 U3016 ( .A(N2590), .B(n2625), .Z(n2679) );
  AO3 U3017 ( .A(n2619), .B(n2681), .C(n2682), .D(n2683), .Z(n3198) );
  AO2 U3018 ( .A(n2623), .B(n448), .C(n4519), .D(n2624), .Z(n2683) );
  ND2 U3019 ( .A(N2591), .B(n2625), .Z(n2682) );
  AO3 U3020 ( .A(n2619), .B(n2684), .C(n2685), .D(n2686), .Z(n3197) );
  AO2 U3021 ( .A(n2623), .B(n447), .C(n4523), .D(n2624), .Z(n2686) );
  ND2 U3022 ( .A(N2592), .B(n2625), .Z(n2685) );
  AO3 U3023 ( .A(n2619), .B(n2687), .C(n2688), .D(n2689), .Z(n3196) );
  AO2 U3024 ( .A(n2623), .B(n446), .C(n4527), .D(n2624), .Z(n2689) );
  ND2 U3025 ( .A(N2593), .B(n2625), .Z(n2688) );
  AO7 U3026 ( .A(n4463), .B(n2690), .C(n2691), .Z(n3195) );
  AO2 U3027 ( .A(n2692), .B(N2579), .C(n2693), .D(n234), .Z(n2691) );
  AO7 U3028 ( .A(n4452), .B(n2690), .C(n2694), .Z(n3194) );
  AO2 U3029 ( .A(n2692), .B(N2580), .C(n2693), .D(n233), .Z(n2694) );
  AO7 U3030 ( .A(n4471), .B(n2690), .C(n2695), .Z(n3193) );
  AO2 U3031 ( .A(n2692), .B(N2581), .C(n2693), .D(n232), .Z(n2695) );
  AO7 U3032 ( .A(n4476), .B(n2690), .C(n2696), .Z(n3192) );
  AO2 U3033 ( .A(n2692), .B(N2582), .C(n2693), .D(n231), .Z(n2696) );
  AO7 U3034 ( .A(n4481), .B(n2690), .C(n2697), .Z(n3191) );
  AO2 U3035 ( .A(n2692), .B(N2583), .C(n2693), .D(n230), .Z(n2697) );
  AO7 U3036 ( .A(n4486), .B(n2690), .C(n2698), .Z(n3190) );
  AO2 U3037 ( .A(n2692), .B(N2584), .C(n2693), .D(n229), .Z(n2698) );
  AO7 U3038 ( .A(n4491), .B(n2690), .C(n2699), .Z(n3189) );
  AO2 U3039 ( .A(n2692), .B(N2585), .C(n2693), .D(n228), .Z(n2699) );
  AO7 U3040 ( .A(n4496), .B(n2690), .C(n2700), .Z(n3188) );
  AO2 U3041 ( .A(n2692), .B(N2586), .C(n2693), .D(n227), .Z(n2700) );
  AO7 U3042 ( .A(n4501), .B(n2690), .C(n2701), .Z(n3187) );
  AO2 U3043 ( .A(n2692), .B(N2587), .C(n2693), .D(n226), .Z(n2701) );
  AO7 U3044 ( .A(n4505), .B(n2690), .C(n2702), .Z(n3186) );
  AO2 U3045 ( .A(n2692), .B(N2588), .C(n2693), .D(n225), .Z(n2702) );
  AO7 U3046 ( .A(n4509), .B(n2690), .C(n2703), .Z(n3185) );
  AO2 U3047 ( .A(n2692), .B(N2589), .C(n2693), .D(n224), .Z(n2703) );
  AO7 U3048 ( .A(n4513), .B(n2690), .C(n2704), .Z(n3184) );
  AO2 U3049 ( .A(n2692), .B(N2590), .C(n2693), .D(n223), .Z(n2704) );
  AO7 U3050 ( .A(n4517), .B(n2690), .C(n2705), .Z(n3183) );
  AO2 U3051 ( .A(n2692), .B(N2591), .C(n2693), .D(n222), .Z(n2705) );
  AO7 U3052 ( .A(n4521), .B(n2690), .C(n2706), .Z(n3182) );
  AO2 U3053 ( .A(n2692), .B(N2592), .C(n2693), .D(n221), .Z(n2706) );
  AO7 U3054 ( .A(n4525), .B(n2690), .C(n2707), .Z(n3181) );
  AO2 U3055 ( .A(n2692), .B(N2593), .C(n2693), .D(n220), .Z(n2707) );
  AO7 U3056 ( .A(n4529), .B(n2690), .C(n2708), .Z(n3180) );
  AO2 U3057 ( .A(n2692), .B(N2594), .C(n2693), .D(n219), .Z(n2708) );
  AO7 U3058 ( .A(n4534), .B(n2690), .C(n2709), .Z(n3179) );
  AO2 U3059 ( .A(N2595), .B(n2692), .C(n2693), .D(n218), .Z(n2709) );
  AO7 U3060 ( .A(n4538), .B(n2690), .C(n2710), .Z(n3178) );
  AO2 U3061 ( .A(N2596), .B(n2692), .C(n2693), .D(n217), .Z(n2710) );
  AO7 U3062 ( .A(n4542), .B(n2690), .C(n2711), .Z(n3177) );
  AO2 U3063 ( .A(N2597), .B(n2692), .C(n2693), .D(n216), .Z(n2711) );
  AO7 U3064 ( .A(n4546), .B(n2690), .C(n2712), .Z(n3176) );
  AO2 U3065 ( .A(N2598), .B(n2692), .C(n2693), .D(n215), .Z(n2712) );
  AO7 U3066 ( .A(n4550), .B(n2690), .C(n2713), .Z(n3175) );
  AO2 U3067 ( .A(N2599), .B(n2692), .C(n2693), .D(n214), .Z(n2713) );
  AO7 U3068 ( .A(n4554), .B(n2690), .C(n2714), .Z(n3174) );
  AO2 U3069 ( .A(N2600), .B(n2692), .C(n2693), .D(n213), .Z(n2714) );
  AO7 U3070 ( .A(n4558), .B(n2690), .C(n2715), .Z(n3173) );
  AO2 U3071 ( .A(N2601), .B(n2692), .C(n2693), .D(n212), .Z(n2715) );
  AO7 U3072 ( .A(n4562), .B(n2690), .C(n2716), .Z(n3172) );
  AO2 U3073 ( .A(N2602), .B(n2692), .C(n2693), .D(n211), .Z(n2716) );
  AO7 U3074 ( .A(n4566), .B(n2690), .C(n2717), .Z(n3171) );
  AO2 U3075 ( .A(N2603), .B(n2692), .C(n2693), .D(n210), .Z(n2717) );
  AO7 U3076 ( .A(n4570), .B(n2690), .C(n2718), .Z(n3170) );
  AO2 U3077 ( .A(N2604), .B(n2692), .C(n2693), .D(n209), .Z(n2718) );
  AO7 U3078 ( .A(n4574), .B(n2690), .C(n2719), .Z(n3169) );
  AO2 U3079 ( .A(N2605), .B(n2692), .C(n2693), .D(n208), .Z(n2719) );
  AO7 U3080 ( .A(n4578), .B(n2690), .C(n2720), .Z(n3168) );
  AO2 U3081 ( .A(N2606), .B(n2692), .C(n2693), .D(n207), .Z(n2720) );
  AO7 U3082 ( .A(n4582), .B(n2690), .C(n2721), .Z(n3167) );
  AO2 U3083 ( .A(N2607), .B(n2692), .C(n2693), .D(n206), .Z(n2721) );
  AO7 U3084 ( .A(n4586), .B(n2690), .C(n2722), .Z(n3166) );
  AO2 U3085 ( .A(N2608), .B(n2692), .C(n2693), .D(n205), .Z(n2722) );
  AO7 U3086 ( .A(n4643), .B(n2690), .C(n2723), .Z(n3165) );
  AO2 U3087 ( .A(N2609), .B(n2692), .C(n2693), .D(n204), .Z(n2723) );
  NR2 U3088 ( .A(n2724), .B(n2725), .Z(n2692) );
  EON1 U3089 ( .A(n4646), .B(n2690), .C(n203), .D(n2693), .Z(n3164) );
  NR2 U3090 ( .A(n2726), .B(n2725), .Z(n2693) );
  IV U3091 ( .A(n2725), .Z(n2690) );
  AO6 U3092 ( .A(n2278), .B(n2254), .C(U3_U21_Z_0), .Z(n2725) );
  AO3 U3093 ( .A(n2619), .B(n2727), .C(n2728), .D(n2729), .Z(n3163) );
  AO2 U3094 ( .A(n2623), .B(n444), .C(n4533), .D(n2624), .Z(n2729) );
  ND2 U3095 ( .A(N2595), .B(n2625), .Z(n2728) );
  AO3 U3096 ( .A(n2619), .B(n2730), .C(n2731), .D(n2732), .Z(n3162) );
  AO2 U3097 ( .A(n2623), .B(n443), .C(n4537), .D(n2624), .Z(n2732) );
  ND2 U3098 ( .A(N2596), .B(n2625), .Z(n2731) );
  AO3 U3099 ( .A(n2619), .B(n2733), .C(n2734), .D(n2735), .Z(n3161) );
  AO2 U3100 ( .A(n2623), .B(n442), .C(n4541), .D(n2624), .Z(n2735) );
  ND2 U3101 ( .A(N2597), .B(n2625), .Z(n2734) );
  AO3 U3102 ( .A(n2619), .B(n2736), .C(n2737), .D(n2738), .Z(n3160) );
  AO2 U3103 ( .A(n2623), .B(n441), .C(n4545), .D(n2624), .Z(n2738) );
  ND2 U3104 ( .A(N2598), .B(n2625), .Z(n2737) );
  AO3 U3105 ( .A(n2619), .B(n2739), .C(n2740), .D(n2741), .Z(n3159) );
  AO2 U3106 ( .A(n2623), .B(n440), .C(n4549), .D(n2624), .Z(n2741) );
  ND2 U3107 ( .A(N2599), .B(n2625), .Z(n2740) );
  AO3 U3108 ( .A(n2619), .B(n2742), .C(n2743), .D(n2744), .Z(n3158) );
  AO2 U3109 ( .A(n2623), .B(n439), .C(n4553), .D(n2624), .Z(n2744) );
  ND2 U3110 ( .A(N2600), .B(n2625), .Z(n2743) );
  AO3 U3111 ( .A(n2619), .B(n2745), .C(n2746), .D(n2747), .Z(n3157) );
  AO2 U3112 ( .A(n2623), .B(n438), .C(n4557), .D(n2624), .Z(n2747) );
  ND2 U3113 ( .A(N2601), .B(n2625), .Z(n2746) );
  AO3 U3114 ( .A(n2619), .B(n2748), .C(n2749), .D(n2750), .Z(n3156) );
  AO2 U3115 ( .A(n2623), .B(n437), .C(n2624), .D(n2205), .Z(n2750) );
  ND2 U3116 ( .A(N2602), .B(n2625), .Z(n2749) );
  IV U3117 ( .A(Datai[23]), .Z(n2748) );
  AO3 U3118 ( .A(n2619), .B(n2751), .C(n2752), .D(n2753), .Z(n3155) );
  AO2 U3119 ( .A(n2623), .B(n436), .C(n2624), .D(n2204), .Z(n2753) );
  ND2 U3120 ( .A(N2603), .B(n2625), .Z(n2752) );
  AO3 U3121 ( .A(n2619), .B(n2754), .C(n2755), .D(n2756), .Z(n3154) );
  AO2 U3122 ( .A(n2623), .B(n435), .C(n2624), .D(n2203), .Z(n2756) );
  ND2 U3123 ( .A(N2604), .B(n2625), .Z(n2755) );
  AO3 U3124 ( .A(n2619), .B(n2757), .C(n2758), .D(n2759), .Z(n3153) );
  AO2 U3125 ( .A(n2623), .B(n434), .C(n2624), .D(n2202), .Z(n2759) );
  ND2 U3126 ( .A(N2605), .B(n2625), .Z(n2758) );
  AO3 U3127 ( .A(n2619), .B(n2760), .C(n2761), .D(n2762), .Z(n3152) );
  AO2 U3128 ( .A(n2623), .B(n433), .C(n2624), .D(n2201), .Z(n2762) );
  ND2 U3129 ( .A(N2606), .B(n2625), .Z(n2761) );
  AO3 U3130 ( .A(n2619), .B(n2763), .C(n2764), .D(n2765), .Z(n3151) );
  AO2 U3131 ( .A(n2623), .B(n432), .C(n2624), .D(n2200), .Z(n2765) );
  ND2 U3132 ( .A(N2607), .B(n2625), .Z(n2764) );
  AO3 U3133 ( .A(n2619), .B(n2766), .C(n2767), .D(n2768), .Z(n3150) );
  AO2 U3134 ( .A(n2623), .B(n431), .C(n2624), .D(n2199), .Z(n2768) );
  ND2 U3135 ( .A(N2608), .B(n2625), .Z(n2767) );
  AO3 U3136 ( .A(n2619), .B(n2769), .C(n2770), .D(n2771), .Z(n3149) );
  AO2 U3137 ( .A(n2623), .B(n430), .C(n2624), .D(n2198), .Z(n2771) );
  ND2 U3138 ( .A(N2609), .B(n2625), .Z(n2770) );
  AO6 U3139 ( .A(n2395), .B(n2772), .C(n2624), .Z(n2625) );
  AO7 U3140 ( .A(n4464), .B(n2773), .C(n2774), .Z(n3148) );
  EO1 U3141 ( .A(n2623), .B(n429), .C(n2775), .D(n2619), .Z(n2774) );
  ND2 U3142 ( .A(n2392), .B(n2773), .Z(n2619) );
  NR2 U3143 ( .A(n2776), .B(n2624), .Z(n2623) );
  IV U3144 ( .A(n2773), .Z(n2624) );
  AO3 U3145 ( .A(n2245), .B(n2772), .C(n2777), .D(n2778), .Z(n2773) );
  ND2 U3146 ( .A(n2278), .B(n2779), .Z(n2777) );
  AO3 U3147 ( .A(n2780), .B(n2781), .C(n2782), .D(n2783), .Z(n3147) );
  AO2 U3148 ( .A(n2784), .B(Datai[0]), .C(N1750), .D(n2785), .Z(n2783) );
  MUX21L U3149 ( .A(n2786), .B(n4413), .S(n2787), .Z(n2782) );
  AO3 U3150 ( .A(n2780), .B(n2788), .C(n2789), .D(n2790), .Z(n3146) );
  AO2 U3151 ( .A(n2784), .B(Datai[1]), .C(N1751), .D(n2785), .Z(n2790) );
  MUX21L U3152 ( .A(n2791), .B(n4425), .S(n2787), .Z(n2789) );
  AO3 U3153 ( .A(n2780), .B(n2792), .C(n2793), .D(n2794), .Z(n3145) );
  AO2 U3154 ( .A(n2784), .B(Datai[2]), .C(N1752), .D(n2785), .Z(n2794) );
  MUX21L U3155 ( .A(n2795), .B(n4664), .S(n2787), .Z(n2793) );
  AO3 U3156 ( .A(n2780), .B(n2796), .C(n2797), .D(n2798), .Z(n3144) );
  AO2 U3157 ( .A(n2784), .B(Datai[3]), .C(N1753), .D(n2785), .Z(n2798) );
  MUX21L U3158 ( .A(n2799), .B(n4663), .S(n2787), .Z(n2797) );
  AO3 U3159 ( .A(n2780), .B(n2800), .C(n2801), .D(n2802), .Z(n3143) );
  AO2 U3160 ( .A(n2784), .B(Datai[4]), .C(N1754), .D(n2785), .Z(n2802) );
  MUX21L U3161 ( .A(n2803), .B(n4662), .S(n2787), .Z(n2801) );
  AO3 U3162 ( .A(n2780), .B(n2804), .C(n2805), .D(n2806), .Z(n3142) );
  AO2 U3163 ( .A(n2784), .B(Datai[5]), .C(N1755), .D(n2785), .Z(n2806) );
  MUX21L U3164 ( .A(n2807), .B(n4661), .S(n2787), .Z(n2805) );
  AO3 U3165 ( .A(n2780), .B(n2808), .C(n2809), .D(n2810), .Z(n3141) );
  AO2 U3166 ( .A(n2784), .B(Datai[6]), .C(N1756), .D(n2785), .Z(n2810) );
  MUX21L U3167 ( .A(n2811), .B(n4660), .S(n2787), .Z(n2809) );
  AO3 U3168 ( .A(n2812), .B(n2780), .C(n2813), .D(n2814), .Z(n3140) );
  AO2 U3169 ( .A(n2784), .B(Datai[7]), .C(n2785), .D(N1757), .Z(n2814) );
  NR4 U3170 ( .A(n2556), .B(n2787), .C(n2815), .D(n2816), .Z(n2784) );
  MUX21L U3171 ( .A(n2271), .B(n4659), .S(n2787), .Z(n2813) );
  NR3 U3172 ( .A(n2817), .B(n2785), .C(n2818), .Z(n2787) );
  AO4 U3173 ( .A(n2819), .B(n2820), .C(n2606), .D(n2821), .Z(n2818) );
  AO3 U3174 ( .A(n2822), .B(n2781), .C(n2823), .D(n2824), .Z(n3139) );
  AO2 U3175 ( .A(n2825), .B(Datai[0]), .C(n2826), .D(N1750), .Z(n2824) );
  MUX21L U3176 ( .A(n2786), .B(n4416), .S(n2827), .Z(n2823) );
  AO3 U3177 ( .A(n2822), .B(n2788), .C(n2828), .D(n2829), .Z(n3138) );
  AO2 U3178 ( .A(n2825), .B(Datai[1]), .C(n2826), .D(N1751), .Z(n2829) );
  MUX21L U3179 ( .A(n2791), .B(n4428), .S(n2827), .Z(n2828) );
  AO3 U3180 ( .A(n2822), .B(n2792), .C(n2830), .D(n2831), .Z(n3137) );
  AO2 U3181 ( .A(n2825), .B(Datai[2]), .C(n2826), .D(N1752), .Z(n2831) );
  MUX21L U3182 ( .A(n2795), .B(n4405), .S(n2827), .Z(n2830) );
  AO3 U3183 ( .A(n2822), .B(n2796), .C(n2832), .D(n2833), .Z(n3136) );
  AO2 U3184 ( .A(n2825), .B(Datai[3]), .C(n2826), .D(N1753), .Z(n2833) );
  MUX21L U3185 ( .A(n2799), .B(n4438), .S(n2827), .Z(n2832) );
  AO3 U3186 ( .A(n2822), .B(n2800), .C(n2834), .D(n2835), .Z(n3135) );
  AO2 U3187 ( .A(n2825), .B(Datai[4]), .C(n2826), .D(N1754), .Z(n2835) );
  MUX21L U3188 ( .A(n2803), .B(n4448), .S(n2827), .Z(n2834) );
  AO3 U3189 ( .A(n2822), .B(n2804), .C(n2836), .D(n2837), .Z(n3134) );
  AO2 U3190 ( .A(n2825), .B(Datai[5]), .C(n2826), .D(N1755), .Z(n2837) );
  MUX21L U3191 ( .A(n2807), .B(n4374), .S(n2827), .Z(n2836) );
  AO3 U3192 ( .A(n2822), .B(n2808), .C(n2838), .D(n2839), .Z(n3133) );
  AO2 U3193 ( .A(n2825), .B(Datai[6]), .C(n2826), .D(N1756), .Z(n2839) );
  MUX21L U3194 ( .A(n2811), .B(n4395), .S(n2827), .Z(n2838) );
  AO3 U3195 ( .A(n2812), .B(n2822), .C(n2840), .D(n2841), .Z(n3132) );
  AO2 U3196 ( .A(n2825), .B(Datai[7]), .C(n2826), .D(N1757), .Z(n2841) );
  NR4 U3197 ( .A(n2556), .B(n2827), .C(n2815), .D(n2842), .Z(n2825) );
  IV U3198 ( .A(n2822), .Z(n2815) );
  MUX21L U3199 ( .A(n2271), .B(n4385), .S(n2827), .Z(n2840) );
  NR3 U3200 ( .A(n2826), .B(n2785), .C(n2843), .Z(n2827) );
  AO4 U3201 ( .A(n2606), .B(n2844), .C(n2819), .D(n2821), .Z(n2843) );
  NR2 U3202 ( .A(n2822), .B(n2590), .Z(n2785) );
  AO3 U3203 ( .A(n2820), .B(n2781), .C(n2845), .D(n2846), .Z(n3131) );
  AO2 U3204 ( .A(n2847), .B(Datai[0]), .C(n2848), .D(N1750), .Z(n2846) );
  MUX21L U3205 ( .A(n2786), .B(n4407), .S(n2849), .Z(n2845) );
  AO3 U3206 ( .A(n2820), .B(n2788), .C(n2850), .D(n2851), .Z(n3130) );
  AO2 U3207 ( .A(n2847), .B(Datai[1]), .C(n2848), .D(N1751), .Z(n2851) );
  MUX21L U3208 ( .A(n2791), .B(n4419), .S(n2849), .Z(n2850) );
  AO3 U3209 ( .A(n2820), .B(n2792), .C(n2852), .D(n2853), .Z(n3129) );
  AO2 U3210 ( .A(n2847), .B(Datai[2]), .C(n2848), .D(N1752), .Z(n2853) );
  MUX21L U3211 ( .A(n2795), .B(n4397), .S(n2849), .Z(n2852) );
  AO3 U3212 ( .A(n2820), .B(n2796), .C(n2854), .D(n2855), .Z(n3128) );
  AO2 U3213 ( .A(n2847), .B(Datai[3]), .C(n2848), .D(N1753), .Z(n2855) );
  MUX21L U3214 ( .A(n2799), .B(n4431), .S(n2849), .Z(n2854) );
  AO3 U3215 ( .A(n2820), .B(n2800), .C(n2856), .D(n2857), .Z(n3127) );
  AO2 U3216 ( .A(n2847), .B(Datai[4]), .C(n2848), .D(N1754), .Z(n2857) );
  MUX21L U3217 ( .A(n2803), .B(n4441), .S(n2849), .Z(n2856) );
  AO3 U3218 ( .A(n2820), .B(n2804), .C(n2858), .D(n2859), .Z(n3126) );
  AO2 U3219 ( .A(n2847), .B(Datai[5]), .C(n2848), .D(N1755), .Z(n2859) );
  MUX21L U3220 ( .A(n2807), .B(n4367), .S(n2849), .Z(n2858) );
  AO3 U3221 ( .A(n2820), .B(n2808), .C(n2860), .D(n2861), .Z(n3125) );
  AO2 U3222 ( .A(n2847), .B(Datai[6]), .C(n2848), .D(N1756), .Z(n2861) );
  MUX21L U3223 ( .A(n2811), .B(n4388), .S(n2849), .Z(n2860) );
  AO3 U3224 ( .A(n2812), .B(n2820), .C(n2862), .D(n2863), .Z(n3124) );
  AO2 U3225 ( .A(n2847), .B(Datai[7]), .C(n2848), .D(N1757), .Z(n2863) );
  NR4 U3226 ( .A(n2556), .B(n2849), .C(n2864), .D(n2842), .Z(n2847) );
  IV U3227 ( .A(n2820), .Z(n2842) );
  MUX21L U3228 ( .A(n2271), .B(n4377), .S(n2849), .Z(n2862) );
  NR3 U3229 ( .A(n2848), .B(n2826), .C(n2865), .Z(n2849) );
  AO4 U3230 ( .A(n2606), .B(n2866), .C(n2819), .D(n2844), .Z(n2865) );
  NR2 U3231 ( .A(n2820), .B(n2590), .Z(n2826) );
  AO3 U3232 ( .A(n2867), .B(n2868), .C(n2869), .D(n2870), .Z(n3123) );
  AO2 U3233 ( .A(n2871), .B(Datai[0]), .C(n2872), .D(n2864), .Z(n2870) );
  MUX21L U3234 ( .A(n2786), .B(n4410), .S(n2873), .Z(n2869) );
  AO3 U3235 ( .A(n2874), .B(n2868), .C(n2875), .D(n2876), .Z(n3122) );
  AO2 U3236 ( .A(n2871), .B(Datai[1]), .C(n2877), .D(n2864), .Z(n2876) );
  MUX21L U3237 ( .A(n2791), .B(n4422), .S(n2873), .Z(n2875) );
  AO3 U3238 ( .A(n2878), .B(n2868), .C(n2879), .D(n2880), .Z(n3121) );
  AO2 U3239 ( .A(n2871), .B(Datai[2]), .C(n2881), .D(n2864), .Z(n2880) );
  MUX21L U3240 ( .A(n2795), .B(n4400), .S(n2873), .Z(n2879) );
  AO3 U3241 ( .A(n2882), .B(n2868), .C(n2883), .D(n2884), .Z(n3120) );
  AO2 U3242 ( .A(n2871), .B(Datai[3]), .C(n2885), .D(n2864), .Z(n2884) );
  MUX21L U3243 ( .A(n2799), .B(n4433), .S(n2873), .Z(n2883) );
  AO3 U3244 ( .A(n2886), .B(n2868), .C(n2887), .D(n2888), .Z(n3119) );
  AO2 U3245 ( .A(n2871), .B(Datai[4]), .C(n2889), .D(n2864), .Z(n2888) );
  MUX21L U3246 ( .A(n2803), .B(n4443), .S(n2873), .Z(n2887) );
  AO3 U3247 ( .A(n2890), .B(n2868), .C(n2891), .D(n2892), .Z(n3118) );
  AO2 U3248 ( .A(n2871), .B(Datai[5]), .C(n2893), .D(n2864), .Z(n2892) );
  MUX21L U3249 ( .A(n2807), .B(n4369), .S(n2873), .Z(n2891) );
  AO3 U3250 ( .A(n2894), .B(n2868), .C(n2895), .D(n2896), .Z(n3117) );
  AO2 U3251 ( .A(n2871), .B(Datai[6]), .C(n2897), .D(n2864), .Z(n2896) );
  MUX21L U3252 ( .A(n2811), .B(n4390), .S(n2873), .Z(n2895) );
  AO3 U3253 ( .A(n2265), .B(n2868), .C(n2898), .D(n2899), .Z(n3116) );
  AO2 U3254 ( .A(n2871), .B(Datai[7]), .C(n2864), .D(n2269), .Z(n2899) );
  NR4 U3255 ( .A(n2556), .B(n2873), .C(n2900), .D(n2864), .Z(n2871) );
  IV U3256 ( .A(n2821), .Z(n2864) );
  MUX21L U3257 ( .A(n2271), .B(n4380), .S(n2873), .Z(n2898) );
  NR3 U3258 ( .A(n2901), .B(n2848), .C(n2902), .Z(n2873) );
  AO4 U3259 ( .A(n2606), .B(n2903), .C(n2819), .D(n2866), .Z(n2902) );
  NR2 U3260 ( .A(n2821), .B(n2590), .Z(n2848) );
  ND2 U3261 ( .A(n2904), .B(n3020), .Z(n2821) );
  AO3 U3262 ( .A(n2867), .B(n3232), .C(n3235), .D(n3237), .Z(n3115) );
  AO2 U3263 ( .A(n3288), .B(Datai[0]), .C(n2900), .D(n2872), .Z(n3237) );
  MUX21L U3264 ( .A(n2786), .B(n4412), .S(n3289), .Z(n3235) );
  AO3 U3265 ( .A(n2874), .B(n3232), .C(n3290), .D(n3291), .Z(n3114) );
  AO2 U3266 ( .A(n3288), .B(Datai[1]), .C(n2900), .D(n2877), .Z(n3291) );
  MUX21L U3267 ( .A(n2791), .B(n4424), .S(n3289), .Z(n3290) );
  AO3 U3268 ( .A(n2878), .B(n3232), .C(n3292), .D(n3293), .Z(n3113) );
  AO2 U3269 ( .A(n3288), .B(Datai[2]), .C(n2900), .D(n2881), .Z(n3293) );
  MUX21L U3270 ( .A(n2795), .B(n4402), .S(n3289), .Z(n3292) );
  AO3 U3271 ( .A(n2882), .B(n3232), .C(n3294), .D(n3295), .Z(n3112) );
  AO2 U3272 ( .A(n3288), .B(Datai[3]), .C(n2900), .D(n2885), .Z(n3295) );
  MUX21L U3273 ( .A(n2799), .B(n4435), .S(n3289), .Z(n3294) );
  AO3 U3274 ( .A(n2886), .B(n3232), .C(n3296), .D(n3297), .Z(n3111) );
  AO2 U3275 ( .A(n3288), .B(Datai[4]), .C(n2900), .D(n2889), .Z(n3297) );
  MUX21L U3276 ( .A(n2803), .B(n4445), .S(n3289), .Z(n3296) );
  AO3 U3277 ( .A(n2890), .B(n3232), .C(n3298), .D(n3299), .Z(n3110) );
  AO2 U3278 ( .A(n3288), .B(Datai[5]), .C(n2900), .D(n2893), .Z(n3299) );
  MUX21L U3279 ( .A(n2807), .B(n4371), .S(n3289), .Z(n3298) );
  AO3 U3280 ( .A(n2894), .B(n3232), .C(n3300), .D(n3301), .Z(n3109) );
  AO2 U3281 ( .A(n3288), .B(Datai[6]), .C(n2900), .D(n2897), .Z(n3301) );
  MUX21L U3282 ( .A(n2811), .B(n4392), .S(n3289), .Z(n3300) );
  AO3 U3283 ( .A(n2265), .B(n3232), .C(n3302), .D(n3303), .Z(n3108) );
  AO2 U3284 ( .A(n3288), .B(Datai[7]), .C(n2900), .D(n2269), .Z(n3303) );
  NR4 U3285 ( .A(n2556), .B(n3289), .C(n3304), .D(n2900), .Z(n3288) );
  MUX21L U3286 ( .A(n2271), .B(n4382), .S(n3289), .Z(n3302) );
  NR3 U3287 ( .A(n3305), .B(n2901), .C(n3306), .Z(n3289) );
  AO4 U3288 ( .A(n2606), .B(n3307), .C(n2819), .D(n2903), .Z(n3306) );
  IV U3289 ( .A(n2868), .Z(n2901) );
  ND2 U3290 ( .A(n2900), .B(n2364), .Z(n2868) );
  IV U3291 ( .A(n2844), .Z(n2900) );
  ND2 U3292 ( .A(n2904), .B(n3308), .Z(n2844) );
  AO3 U3293 ( .A(n2867), .B(n3309), .C(n3310), .D(n3311), .Z(n3107) );
  AO2 U3294 ( .A(n3312), .B(Datai[0]), .C(n3304), .D(n2872), .Z(n3311) );
  MUX21L U3295 ( .A(n2786), .B(n4594), .S(n3313), .Z(n3310) );
  AO3 U3296 ( .A(n2874), .B(n3309), .C(n3314), .D(n3315), .Z(n3106) );
  AO2 U3297 ( .A(n3312), .B(Datai[1]), .C(n3304), .D(n2877), .Z(n3315) );
  MUX21L U3298 ( .A(n2791), .B(n4599), .S(n3313), .Z(n3314) );
  AO3 U3299 ( .A(n2878), .B(n3309), .C(n3316), .D(n3317), .Z(n3105) );
  AO2 U3300 ( .A(n3312), .B(Datai[2]), .C(n3304), .D(n2881), .Z(n3317) );
  MUX21L U3301 ( .A(n2795), .B(n4605), .S(n3313), .Z(n3316) );
  AO3 U3302 ( .A(n2882), .B(n3309), .C(n3318), .D(n3319), .Z(n3104) );
  AO2 U3303 ( .A(n3312), .B(Datai[3]), .C(n3304), .D(n2885), .Z(n3319) );
  MUX21L U3304 ( .A(n2799), .B(n4611), .S(n3313), .Z(n3318) );
  AO3 U3305 ( .A(n2886), .B(n3309), .C(n3320), .D(n3321), .Z(n3103) );
  AO2 U3306 ( .A(n3312), .B(Datai[4]), .C(n3304), .D(n2889), .Z(n3321) );
  MUX21L U3307 ( .A(n2803), .B(n4617), .S(n3313), .Z(n3320) );
  AO3 U3308 ( .A(n2890), .B(n3309), .C(n3322), .D(n3323), .Z(n3102) );
  AO2 U3309 ( .A(n3312), .B(Datai[5]), .C(n3304), .D(n2893), .Z(n3323) );
  MUX21L U3310 ( .A(n2807), .B(n4623), .S(n3313), .Z(n3322) );
  AO3 U3311 ( .A(n2894), .B(n3309), .C(n3324), .D(n3325), .Z(n3101) );
  AO2 U3312 ( .A(n3312), .B(Datai[6]), .C(n3304), .D(n2897), .Z(n3325) );
  MUX21L U3313 ( .A(n2811), .B(n4630), .S(n3313), .Z(n3324) );
  AO3 U3314 ( .A(n2265), .B(n3309), .C(n3326), .D(n3327), .Z(n3100) );
  AO2 U3315 ( .A(n3312), .B(Datai[7]), .C(n3304), .D(n2269), .Z(n3327) );
  NR4 U3316 ( .A(n2556), .B(n3313), .C(n3328), .D(n3304), .Z(n3312) );
  MUX21L U3317 ( .A(n2271), .B(n4635), .S(n3313), .Z(n3326) );
  NR3 U3318 ( .A(n3329), .B(n3305), .C(n3330), .Z(n3313) );
  AO4 U3319 ( .A(n2606), .B(n3331), .C(n2819), .D(n3307), .Z(n3330) );
  IV U3320 ( .A(n3232), .Z(n3305) );
  ND2 U3321 ( .A(n3304), .B(n2364), .Z(n3232) );
  IV U3322 ( .A(n2866), .Z(n3304) );
  ND2 U3323 ( .A(n2904), .B(n3332), .Z(n2866) );
  AO3 U3324 ( .A(n2867), .B(n3333), .C(n3334), .D(n3335), .Z(n3099) );
  AO2 U3325 ( .A(n3336), .B(Datai[0]), .C(n3328), .D(n2872), .Z(n3335) );
  MUX21L U3326 ( .A(n2786), .B(n4593), .S(n3337), .Z(n3334) );
  AO3 U3327 ( .A(n2874), .B(n3333), .C(n3338), .D(n3339), .Z(n3098) );
  AO2 U3328 ( .A(n3336), .B(Datai[1]), .C(n3328), .D(n2877), .Z(n3339) );
  MUX21L U3329 ( .A(n2791), .B(n4598), .S(n3337), .Z(n3338) );
  AO3 U3330 ( .A(n2878), .B(n3333), .C(n3340), .D(n3341), .Z(n3097) );
  AO2 U3331 ( .A(n3336), .B(Datai[2]), .C(n3328), .D(n2881), .Z(n3341) );
  MUX21L U3332 ( .A(n2795), .B(n4604), .S(n3337), .Z(n3340) );
  AO3 U3333 ( .A(n2882), .B(n3333), .C(n3342), .D(n3343), .Z(n3096) );
  AO2 U3334 ( .A(n3336), .B(Datai[3]), .C(n3328), .D(n2885), .Z(n3343) );
  MUX21L U3335 ( .A(n2799), .B(n4610), .S(n3337), .Z(n3342) );
  AO3 U3336 ( .A(n2886), .B(n3333), .C(n3344), .D(n3345), .Z(n3095) );
  AO2 U3337 ( .A(n3336), .B(Datai[4]), .C(n3328), .D(n2889), .Z(n3345) );
  MUX21L U3338 ( .A(n2803), .B(n4616), .S(n3337), .Z(n3344) );
  AO3 U3339 ( .A(n2890), .B(n3333), .C(n3346), .D(n3347), .Z(n3094) );
  AO2 U3340 ( .A(n3336), .B(Datai[5]), .C(n3328), .D(n2893), .Z(n3347) );
  MUX21L U3341 ( .A(n2807), .B(n4622), .S(n3337), .Z(n3346) );
  AO3 U3342 ( .A(n2894), .B(n3333), .C(n3348), .D(n3349), .Z(n3093) );
  AO2 U3343 ( .A(n3336), .B(Datai[6]), .C(n3328), .D(n2897), .Z(n3349) );
  MUX21L U3344 ( .A(n2811), .B(n4629), .S(n3337), .Z(n3348) );
  AO3 U3345 ( .A(n2265), .B(n3333), .C(n3350), .D(n3351), .Z(n3092) );
  AO2 U3346 ( .A(n3336), .B(Datai[7]), .C(n3328), .D(n2269), .Z(n3351) );
  NR4 U3347 ( .A(n2556), .B(n3337), .C(n3352), .D(n3328), .Z(n3336) );
  MUX21L U3348 ( .A(n2271), .B(n4634), .S(n3337), .Z(n3350) );
  NR3 U3349 ( .A(n3353), .B(n3329), .C(n3354), .Z(n3337) );
  AO4 U3350 ( .A(n2606), .B(n3355), .C(n2819), .D(n3331), .Z(n3354) );
  IV U3351 ( .A(n3309), .Z(n3329) );
  ND2 U3352 ( .A(n3328), .B(n2364), .Z(n3309) );
  IV U3353 ( .A(n2903), .Z(n3328) );
  ND2 U3354 ( .A(n2904), .B(n3356), .Z(n2903) );
  NR2 U3355 ( .A(n2171), .B(n2147), .Z(n2904) );
  AO3 U3356 ( .A(n2867), .B(n3357), .C(n3358), .D(n3359), .Z(n3091) );
  AO2 U3357 ( .A(n3360), .B(Datai[0]), .C(n3352), .D(n2872), .Z(n3359) );
  MUX21L U3358 ( .A(n2786), .B(n4592), .S(n3361), .Z(n3358) );
  AO3 U3359 ( .A(n2874), .B(n3357), .C(n3362), .D(n3363), .Z(n3090) );
  AO2 U3360 ( .A(n3360), .B(Datai[1]), .C(n3352), .D(n2877), .Z(n3363) );
  MUX21L U3361 ( .A(n2791), .B(n4597), .S(n3361), .Z(n3362) );
  AO3 U3362 ( .A(n2878), .B(n3357), .C(n3364), .D(n3365), .Z(n3089) );
  AO2 U3363 ( .A(n3360), .B(Datai[2]), .C(n3352), .D(n2881), .Z(n3365) );
  MUX21L U3364 ( .A(n2795), .B(n4603), .S(n3361), .Z(n3364) );
  AO3 U3365 ( .A(n2882), .B(n3357), .C(n3366), .D(n3367), .Z(n3088) );
  AO2 U3366 ( .A(n3360), .B(Datai[3]), .C(n3352), .D(n2885), .Z(n3367) );
  MUX21L U3367 ( .A(n2799), .B(n4609), .S(n3361), .Z(n3366) );
  AO3 U3368 ( .A(n2886), .B(n3357), .C(n3368), .D(n3369), .Z(n3087) );
  AO2 U3369 ( .A(n3360), .B(Datai[4]), .C(n3352), .D(n2889), .Z(n3369) );
  MUX21L U3370 ( .A(n2803), .B(n4615), .S(n3361), .Z(n3368) );
  AO3 U3371 ( .A(n2890), .B(n3357), .C(n3370), .D(n3371), .Z(n3086) );
  AO2 U3372 ( .A(n3360), .B(Datai[5]), .C(n3352), .D(n2893), .Z(n3371) );
  MUX21L U3373 ( .A(n2807), .B(n4621), .S(n3361), .Z(n3370) );
  AO3 U3374 ( .A(n2894), .B(n3357), .C(n3372), .D(n3373), .Z(n3085) );
  AO2 U3375 ( .A(n3360), .B(Datai[6]), .C(n3352), .D(n2897), .Z(n3373) );
  MUX21L U3376 ( .A(n2811), .B(n4628), .S(n3361), .Z(n3372) );
  AO3 U3377 ( .A(n2265), .B(n3357), .C(n3374), .D(n3375), .Z(n3084) );
  AO2 U3378 ( .A(n3360), .B(Datai[7]), .C(n3352), .D(n2269), .Z(n3375) );
  NR4 U3379 ( .A(n2556), .B(n3361), .C(n3376), .D(n3352), .Z(n3360) );
  MUX21L U3380 ( .A(n2271), .B(n4633), .S(n3361), .Z(n3374) );
  NR3 U3381 ( .A(n3377), .B(n3353), .C(n3378), .Z(n3361) );
  AO4 U3382 ( .A(n2606), .B(n3379), .C(n2819), .D(n3355), .Z(n3378) );
  IV U3383 ( .A(n3333), .Z(n3353) );
  ND2 U3384 ( .A(n3352), .B(n2364), .Z(n3333) );
  IV U3385 ( .A(n3307), .Z(n3352) );
  ND2 U3386 ( .A(n3380), .B(n3020), .Z(n3307) );
  AO3 U3387 ( .A(n2867), .B(n3381), .C(n3382), .D(n3383), .Z(n3083) );
  AO2 U3388 ( .A(n3384), .B(Datai[0]), .C(n3376), .D(n2872), .Z(n3383) );
  MUX21L U3389 ( .A(n2786), .B(n4591), .S(n3385), .Z(n3382) );
  AO3 U3390 ( .A(n2874), .B(n3381), .C(n3386), .D(n3387), .Z(n3082) );
  AO2 U3391 ( .A(n3384), .B(Datai[1]), .C(n3376), .D(n2877), .Z(n3387) );
  MUX21L U3392 ( .A(n2791), .B(n4596), .S(n3385), .Z(n3386) );
  AO3 U3393 ( .A(n2878), .B(n3381), .C(n3388), .D(n3389), .Z(n3081) );
  AO2 U3394 ( .A(n3384), .B(Datai[2]), .C(n3376), .D(n2881), .Z(n3389) );
  MUX21L U3395 ( .A(n2795), .B(n4602), .S(n3385), .Z(n3388) );
  AO3 U3396 ( .A(n2882), .B(n3381), .C(n3390), .D(n3391), .Z(n3080) );
  AO2 U3397 ( .A(n3384), .B(Datai[3]), .C(n3376), .D(n2885), .Z(n3391) );
  MUX21L U3398 ( .A(n2799), .B(n4608), .S(n3385), .Z(n3390) );
  AO3 U3399 ( .A(n2886), .B(n3381), .C(n3392), .D(n3393), .Z(n3079) );
  AO2 U3400 ( .A(n3384), .B(Datai[4]), .C(n3376), .D(n2889), .Z(n3393) );
  MUX21L U3401 ( .A(n2803), .B(n4614), .S(n3385), .Z(n3392) );
  AO3 U3402 ( .A(n2890), .B(n3381), .C(n3394), .D(n3395), .Z(n3078) );
  AO2 U3403 ( .A(n3384), .B(Datai[5]), .C(n3376), .D(n2893), .Z(n3395) );
  MUX21L U3404 ( .A(n2807), .B(n4620), .S(n3385), .Z(n3394) );
  AO3 U3405 ( .A(n2894), .B(n3381), .C(n3396), .D(n3397), .Z(n3077) );
  AO2 U3406 ( .A(n3384), .B(Datai[6]), .C(n3376), .D(n2897), .Z(n3397) );
  MUX21L U3407 ( .A(n2811), .B(n4627), .S(n3385), .Z(n3396) );
  AO3 U3408 ( .A(n2265), .B(n3381), .C(n3398), .D(n3399), .Z(n3076) );
  AO2 U3409 ( .A(n3384), .B(Datai[7]), .C(n3376), .D(n2269), .Z(n3399) );
  NR4 U3410 ( .A(n2556), .B(n3385), .C(n3400), .D(n3376), .Z(n3384) );
  MUX21L U3411 ( .A(n2271), .B(n4632), .S(n3385), .Z(n3398) );
  NR3 U3412 ( .A(n3401), .B(n3377), .C(n3402), .Z(n3385) );
  AO4 U3413 ( .A(n2606), .B(n3403), .C(n2819), .D(n3379), .Z(n3402) );
  IV U3414 ( .A(n3357), .Z(n3377) );
  ND2 U3415 ( .A(n3376), .B(n2364), .Z(n3357) );
  IV U3416 ( .A(n3331), .Z(n3376) );
  ND2 U3417 ( .A(n3380), .B(n3308), .Z(n3331) );
  AO3 U3418 ( .A(n2867), .B(n3404), .C(n3405), .D(n3406), .Z(n3075) );
  AO2 U3419 ( .A(n3407), .B(Datai[0]), .C(n3400), .D(n2872), .Z(n3406) );
  MUX21L U3420 ( .A(n2786), .B(n4417), .S(n3408), .Z(n3405) );
  AO3 U3421 ( .A(n2874), .B(n3404), .C(n3409), .D(n3410), .Z(n3074) );
  AO2 U3422 ( .A(n3407), .B(Datai[1]), .C(n3400), .D(n2877), .Z(n3410) );
  MUX21L U3423 ( .A(n2791), .B(n4429), .S(n3408), .Z(n3409) );
  AO3 U3424 ( .A(n2878), .B(n3404), .C(n3411), .D(n3412), .Z(n3073) );
  AO2 U3425 ( .A(n3407), .B(Datai[2]), .C(n3400), .D(n2881), .Z(n3412) );
  MUX21L U3426 ( .A(n2795), .B(n4601), .S(n3408), .Z(n3411) );
  AO3 U3427 ( .A(n2882), .B(n3404), .C(n3413), .D(n3414), .Z(n3072) );
  AO2 U3428 ( .A(n3407), .B(Datai[3]), .C(n3400), .D(n2885), .Z(n3414) );
  MUX21L U3429 ( .A(n2799), .B(n4439), .S(n3408), .Z(n3413) );
  AO3 U3430 ( .A(n2886), .B(n3404), .C(n3415), .D(n3416), .Z(n3071) );
  AO2 U3431 ( .A(n3407), .B(Datai[4]), .C(n3400), .D(n2889), .Z(n3416) );
  MUX21L U3432 ( .A(n2803), .B(n4449), .S(n3408), .Z(n3415) );
  AO3 U3433 ( .A(n2890), .B(n3404), .C(n3417), .D(n3418), .Z(n3070) );
  AO2 U3434 ( .A(n3407), .B(Datai[5]), .C(n3400), .D(n2893), .Z(n3418) );
  MUX21L U3435 ( .A(n2807), .B(n4375), .S(n3408), .Z(n3417) );
  AO3 U3436 ( .A(n2894), .B(n3404), .C(n3419), .D(n3420), .Z(n3069) );
  AO2 U3437 ( .A(n3407), .B(Datai[6]), .C(n3400), .D(n2897), .Z(n3420) );
  MUX21L U3438 ( .A(n2811), .B(n4626), .S(n3408), .Z(n3419) );
  AO3 U3439 ( .A(n2265), .B(n3404), .C(n3421), .D(n3422), .Z(n3068) );
  AO2 U3440 ( .A(n3407), .B(Datai[7]), .C(n3400), .D(n2269), .Z(n3422) );
  NR4 U3441 ( .A(n2556), .B(n3408), .C(n3423), .D(n3400), .Z(n3407) );
  MUX21L U3442 ( .A(n2271), .B(n4386), .S(n3408), .Z(n3421) );
  NR3 U3443 ( .A(n3424), .B(n3401), .C(n3425), .Z(n3408) );
  AO4 U3444 ( .A(n2606), .B(n3426), .C(n2819), .D(n3403), .Z(n3425) );
  IV U3445 ( .A(n3381), .Z(n3401) );
  ND2 U3446 ( .A(n3400), .B(n2364), .Z(n3381) );
  IV U3447 ( .A(n3355), .Z(n3400) );
  ND2 U3448 ( .A(n3380), .B(n3332), .Z(n3355) );
  AO3 U3449 ( .A(n2867), .B(n3427), .C(n3428), .D(n3429), .Z(n3067) );
  AO2 U3450 ( .A(n3430), .B(Datai[0]), .C(n3423), .D(n2872), .Z(n3429) );
  MUX21L U3451 ( .A(n2786), .B(n4408), .S(n3431), .Z(n3428) );
  AO3 U3452 ( .A(n2874), .B(n3427), .C(n3432), .D(n3433), .Z(n3066) );
  AO2 U3453 ( .A(n3430), .B(Datai[1]), .C(n3423), .D(n2877), .Z(n3433) );
  MUX21L U3454 ( .A(n2791), .B(n4420), .S(n3431), .Z(n3432) );
  AO3 U3455 ( .A(n2878), .B(n3427), .C(n3434), .D(n3435), .Z(n3065) );
  AO2 U3456 ( .A(n3430), .B(Datai[2]), .C(n3423), .D(n2881), .Z(n3435) );
  MUX21L U3457 ( .A(n2795), .B(n4398), .S(n3431), .Z(n3434) );
  AO3 U3458 ( .A(n2882), .B(n3427), .C(n3436), .D(n3437), .Z(n3064) );
  AO2 U3459 ( .A(n3430), .B(Datai[3]), .C(n3423), .D(n2885), .Z(n3437) );
  MUX21L U3460 ( .A(n2799), .B(n4607), .S(n3431), .Z(n3436) );
  AO3 U3461 ( .A(n2886), .B(n3427), .C(n3438), .D(n3439), .Z(n3063) );
  AO2 U3462 ( .A(n3430), .B(Datai[4]), .C(n3423), .D(n2889), .Z(n3439) );
  MUX21L U3463 ( .A(n2803), .B(n4613), .S(n3431), .Z(n3438) );
  AO3 U3464 ( .A(n2890), .B(n3427), .C(n3440), .D(n3441), .Z(n3062) );
  AO2 U3465 ( .A(n3430), .B(Datai[5]), .C(n3423), .D(n2893), .Z(n3441) );
  MUX21L U3466 ( .A(n2807), .B(n4619), .S(n3431), .Z(n3440) );
  AO3 U3467 ( .A(n2894), .B(n3427), .C(n3442), .D(n3443), .Z(n3061) );
  AO2 U3468 ( .A(n3430), .B(Datai[6]), .C(n3423), .D(n2897), .Z(n3443) );
  MUX21L U3469 ( .A(n2811), .B(n4625), .S(n3431), .Z(n3442) );
  AO3 U3470 ( .A(n2265), .B(n3427), .C(n3444), .D(n3445), .Z(n3060) );
  AO2 U3471 ( .A(n3430), .B(Datai[7]), .C(n3423), .D(n2269), .Z(n3445) );
  NR4 U3472 ( .A(n2556), .B(n3431), .C(n3446), .D(n3423), .Z(n3430) );
  MUX21L U3473 ( .A(n2271), .B(n4378), .S(n3431), .Z(n3444) );
  NR3 U3474 ( .A(n3447), .B(n3424), .C(n3448), .Z(n3431) );
  AO4 U3475 ( .A(n2606), .B(n3449), .C(n2819), .D(n3426), .Z(n3448) );
  IV U3476 ( .A(n3404), .Z(n3424) );
  ND2 U3477 ( .A(n3423), .B(n2364), .Z(n3404) );
  IV U3478 ( .A(n3379), .Z(n3423) );
  ND2 U3479 ( .A(n3380), .B(n3356), .Z(n3379) );
  IV U3480 ( .A(n2602), .Z(n3380) );
  ND2 U3481 ( .A(n4457), .B(n2147), .Z(n2602) );
  AO3 U3482 ( .A(n2867), .B(n3450), .C(n3451), .D(n3452), .Z(n3059) );
  AO2 U3483 ( .A(n3453), .B(Datai[0]), .C(n3446), .D(n2872), .Z(n3452) );
  MUX21L U3484 ( .A(n2786), .B(n4411), .S(n3454), .Z(n3451) );
  AO3 U3485 ( .A(n2874), .B(n3450), .C(n3455), .D(n3456), .Z(n3058) );
  AO2 U3486 ( .A(n3453), .B(Datai[1]), .C(n3446), .D(n2877), .Z(n3456) );
  MUX21L U3487 ( .A(n2791), .B(n4423), .S(n3454), .Z(n3455) );
  AO3 U3488 ( .A(n2878), .B(n3450), .C(n3457), .D(n3458), .Z(n3057) );
  AO2 U3489 ( .A(n3453), .B(Datai[2]), .C(n3446), .D(n2881), .Z(n3458) );
  MUX21L U3490 ( .A(n2795), .B(n4401), .S(n3454), .Z(n3457) );
  AO3 U3491 ( .A(n2882), .B(n3450), .C(n3459), .D(n3460), .Z(n3056) );
  AO2 U3492 ( .A(n3453), .B(Datai[3]), .C(n3446), .D(n2885), .Z(n3460) );
  MUX21L U3493 ( .A(n2799), .B(n4434), .S(n3454), .Z(n3459) );
  AO3 U3494 ( .A(n2886), .B(n3450), .C(n3461), .D(n3462), .Z(n3055) );
  AO2 U3495 ( .A(n3453), .B(Datai[4]), .C(n3446), .D(n2889), .Z(n3462) );
  MUX21L U3496 ( .A(n2803), .B(n4444), .S(n3454), .Z(n3461) );
  AO3 U3497 ( .A(n2890), .B(n3450), .C(n3463), .D(n3464), .Z(n3054) );
  AO2 U3498 ( .A(n3453), .B(Datai[5]), .C(n3446), .D(n2893), .Z(n3464) );
  MUX21L U3499 ( .A(n2807), .B(n4370), .S(n3454), .Z(n3463) );
  AO3 U3500 ( .A(n2894), .B(n3450), .C(n3465), .D(n3466), .Z(n3053) );
  AO2 U3501 ( .A(n3453), .B(Datai[6]), .C(n3446), .D(n2897), .Z(n3466) );
  MUX21L U3502 ( .A(n2811), .B(n4391), .S(n3454), .Z(n3465) );
  AO3 U3503 ( .A(n2265), .B(n3450), .C(n3467), .D(n3468), .Z(n3052) );
  AO2 U3504 ( .A(n3453), .B(Datai[7]), .C(n3446), .D(n2269), .Z(n3468) );
  NR4 U3505 ( .A(n2556), .B(n3454), .C(n3469), .D(n3446), .Z(n3453) );
  MUX21L U3506 ( .A(n2271), .B(n4381), .S(n3454), .Z(n3467) );
  NR3 U3507 ( .A(n3470), .B(n3447), .C(n3471), .Z(n3454) );
  AO4 U3508 ( .A(n2606), .B(n3472), .C(n2819), .D(n3449), .Z(n3471) );
  IV U3509 ( .A(n3427), .Z(n3447) );
  ND2 U3510 ( .A(n3446), .B(n2364), .Z(n3427) );
  IV U3511 ( .A(n3403), .Z(n3446) );
  ND2 U3512 ( .A(n3473), .B(n3020), .Z(n3403) );
  AO3 U3513 ( .A(n2867), .B(n3474), .C(n3475), .D(n3476), .Z(n3051) );
  AO2 U3514 ( .A(n3477), .B(Datai[0]), .C(n3469), .D(n2872), .Z(n3476) );
  MUX21L U3515 ( .A(n2786), .B(n4414), .S(n3478), .Z(n3475) );
  AO3 U3516 ( .A(n2874), .B(n3474), .C(n3479), .D(n3480), .Z(n3050) );
  AO2 U3517 ( .A(n3477), .B(Datai[1]), .C(n3469), .D(n2877), .Z(n3480) );
  MUX21L U3518 ( .A(n2791), .B(n4426), .S(n3478), .Z(n3479) );
  AO3 U3519 ( .A(n2878), .B(n3474), .C(n3481), .D(n3482), .Z(n3049) );
  AO2 U3520 ( .A(n3477), .B(Datai[2]), .C(n3469), .D(n2881), .Z(n3482) );
  MUX21L U3521 ( .A(n2795), .B(n4403), .S(n3478), .Z(n3481) );
  AO3 U3522 ( .A(n2882), .B(n3474), .C(n3483), .D(n3484), .Z(n3048) );
  AO2 U3523 ( .A(n3477), .B(Datai[3]), .C(n3469), .D(n2885), .Z(n3484) );
  MUX21L U3524 ( .A(n2799), .B(n4436), .S(n3478), .Z(n3483) );
  AO3 U3525 ( .A(n2886), .B(n3474), .C(n3485), .D(n3486), .Z(n3047) );
  AO2 U3526 ( .A(n3477), .B(Datai[4]), .C(n3469), .D(n2889), .Z(n3486) );
  MUX21L U3527 ( .A(n2803), .B(n4446), .S(n3478), .Z(n3485) );
  AO3 U3528 ( .A(n2890), .B(n3474), .C(n3487), .D(n3488), .Z(n3046) );
  AO2 U3529 ( .A(n3477), .B(Datai[5]), .C(n3469), .D(n2893), .Z(n3488) );
  MUX21L U3530 ( .A(n2807), .B(n4372), .S(n3478), .Z(n3487) );
  AO3 U3531 ( .A(n2894), .B(n3474), .C(n3489), .D(n3490), .Z(n3045) );
  AO2 U3532 ( .A(n3477), .B(Datai[6]), .C(n3469), .D(n2897), .Z(n3490) );
  MUX21L U3533 ( .A(n2811), .B(n4393), .S(n3478), .Z(n3489) );
  AO3 U3534 ( .A(n2265), .B(n3474), .C(n3491), .D(n3492), .Z(n3044) );
  AO2 U3535 ( .A(n3477), .B(Datai[7]), .C(n3469), .D(n2269), .Z(n3492) );
  NR4 U3536 ( .A(n2556), .B(n3478), .C(n3493), .D(n3469), .Z(n3477) );
  MUX21L U3537 ( .A(n2271), .B(n4383), .S(n3478), .Z(n3491) );
  NR3 U3538 ( .A(n3494), .B(n3470), .C(n3495), .Z(n3478) );
  AO4 U3539 ( .A(n2606), .B(n3496), .C(n2819), .D(n3472), .Z(n3495) );
  IV U3540 ( .A(n3450), .Z(n3470) );
  ND2 U3541 ( .A(n3469), .B(n2364), .Z(n3450) );
  IV U3542 ( .A(n3426), .Z(n3469) );
  ND2 U3543 ( .A(n3473), .B(n3308), .Z(n3426) );
  AO3 U3544 ( .A(n2867), .B(n3497), .C(n3498), .D(n3499), .Z(n3043) );
  AO2 U3545 ( .A(n3500), .B(Datai[0]), .C(n3493), .D(n2872), .Z(n3499) );
  MUX21L U3546 ( .A(n2786), .B(n4415), .S(n3501), .Z(n3498) );
  AO3 U3547 ( .A(n2874), .B(n3497), .C(n3502), .D(n3503), .Z(n3042) );
  AO2 U3548 ( .A(n3500), .B(Datai[1]), .C(n3493), .D(n2877), .Z(n3503) );
  MUX21L U3549 ( .A(n2791), .B(n4427), .S(n3501), .Z(n3502) );
  AO3 U3550 ( .A(n2878), .B(n3497), .C(n3504), .D(n3505), .Z(n3041) );
  AO2 U3551 ( .A(n3500), .B(Datai[2]), .C(n3493), .D(n2881), .Z(n3505) );
  MUX21L U3552 ( .A(n2795), .B(n4404), .S(n3501), .Z(n3504) );
  AO3 U3553 ( .A(n2882), .B(n3497), .C(n3506), .D(n3507), .Z(n3040) );
  AO2 U3554 ( .A(n3500), .B(Datai[3]), .C(n3493), .D(n2885), .Z(n3507) );
  MUX21L U3555 ( .A(n2799), .B(n4437), .S(n3501), .Z(n3506) );
  AO3 U3556 ( .A(n2886), .B(n3497), .C(n3508), .D(n3509), .Z(n3039) );
  AO2 U3557 ( .A(n3500), .B(Datai[4]), .C(n3493), .D(n2889), .Z(n3509) );
  MUX21L U3558 ( .A(n2803), .B(n4447), .S(n3501), .Z(n3508) );
  AO3 U3559 ( .A(n2890), .B(n3497), .C(n3510), .D(n3511), .Z(n3038) );
  AO2 U3560 ( .A(n3500), .B(Datai[5]), .C(n3493), .D(n2893), .Z(n3511) );
  MUX21L U3561 ( .A(n2807), .B(n4373), .S(n3501), .Z(n3510) );
  AO3 U3562 ( .A(n2894), .B(n3497), .C(n3512), .D(n3513), .Z(n3037) );
  AO2 U3563 ( .A(n3500), .B(Datai[6]), .C(n3493), .D(n2897), .Z(n3513) );
  MUX21L U3564 ( .A(n2811), .B(n4394), .S(n3501), .Z(n3512) );
  AO3 U3565 ( .A(n2265), .B(n3497), .C(n3514), .D(n3515), .Z(n3036) );
  AO2 U3566 ( .A(n3500), .B(Datai[7]), .C(n3493), .D(n2269), .Z(n3515) );
  NR4 U3567 ( .A(n2556), .B(n3501), .C(n3516), .D(n3493), .Z(n3500) );
  MUX21L U3568 ( .A(n2271), .B(n4384), .S(n3501), .Z(n3514) );
  NR3 U3569 ( .A(n3517), .B(n3494), .C(n3518), .Z(n3501) );
  AO4 U3570 ( .A(n2819), .B(n3496), .C(n2606), .D(n2780), .Z(n3518) );
  IV U3571 ( .A(n3474), .Z(n3494) );
  ND2 U3572 ( .A(n3493), .B(n2364), .Z(n3474) );
  IV U3573 ( .A(n3449), .Z(n3493) );
  ND2 U3574 ( .A(n3473), .B(n3332), .Z(n3449) );
  AO3 U3575 ( .A(n2867), .B(n3519), .C(n3520), .D(n3521), .Z(n3035) );
  AO2 U3576 ( .A(n3522), .B(Datai[0]), .C(n3516), .D(n2872), .Z(n3521) );
  MUX21L U3577 ( .A(n2786), .B(n4406), .S(n3523), .Z(n3520) );
  AO3 U3578 ( .A(n2874), .B(n3519), .C(n3524), .D(n3525), .Z(n3034) );
  AO2 U3579 ( .A(n3522), .B(Datai[1]), .C(n3516), .D(n2877), .Z(n3525) );
  MUX21L U3580 ( .A(n2791), .B(n4418), .S(n3523), .Z(n3524) );
  AO3 U3581 ( .A(n2878), .B(n3519), .C(n3526), .D(n3527), .Z(n3033) );
  AO2 U3582 ( .A(n3522), .B(Datai[2]), .C(n3516), .D(n2881), .Z(n3527) );
  MUX21L U3583 ( .A(n2795), .B(n4396), .S(n3523), .Z(n3526) );
  AO3 U3584 ( .A(n2882), .B(n3519), .C(n3528), .D(n3529), .Z(n3032) );
  AO2 U3585 ( .A(n3522), .B(Datai[3]), .C(n3516), .D(n2885), .Z(n3529) );
  MUX21L U3586 ( .A(n2799), .B(n4430), .S(n3523), .Z(n3528) );
  AO3 U3587 ( .A(n2886), .B(n3519), .C(n3530), .D(n3531), .Z(n3031) );
  AO2 U3588 ( .A(n3522), .B(Datai[4]), .C(n3516), .D(n2889), .Z(n3531) );
  MUX21L U3589 ( .A(n2803), .B(n4440), .S(n3523), .Z(n3530) );
  AO3 U3590 ( .A(n2890), .B(n3519), .C(n3532), .D(n3533), .Z(n3030) );
  AO2 U3591 ( .A(n3522), .B(Datai[5]), .C(n3516), .D(n2893), .Z(n3533) );
  MUX21L U3592 ( .A(n2807), .B(n4366), .S(n3523), .Z(n3532) );
  AO3 U3593 ( .A(n2894), .B(n3519), .C(n3534), .D(n3535), .Z(n3029) );
  AO2 U3594 ( .A(n3522), .B(Datai[6]), .C(n3516), .D(n2897), .Z(n3535) );
  MUX21L U3595 ( .A(n2811), .B(n4387), .S(n3523), .Z(n3534) );
  AO3 U3596 ( .A(n2265), .B(n3519), .C(n3536), .D(n3537), .Z(n3028) );
  AO2 U3597 ( .A(n3516), .B(n2269), .C(n3522), .D(Datai[7]), .Z(n3537) );
  NR4 U3598 ( .A(n2556), .B(n3523), .C(n3516), .D(n2268), .Z(n3522) );
  IV U3599 ( .A(n2812), .Z(n2269) );
  ND2 U3600 ( .A(N819), .B(n2364), .Z(n2812) );
  MUX21L U3601 ( .A(n2271), .B(n4376), .S(n3523), .Z(n3536) );
  NR3 U3602 ( .A(n3538), .B(n3517), .C(n3539), .Z(n3523) );
  AO4 U3603 ( .A(n2819), .B(n2780), .C(n2606), .D(n2822), .Z(n3539) );
  IV U3604 ( .A(n3497), .Z(n3517) );
  ND2 U3605 ( .A(n3516), .B(n2364), .Z(n3497) );
  IV U3606 ( .A(n3472), .Z(n3516) );
  ND2 U3607 ( .A(n3473), .B(n3356), .Z(n3472) );
  NR2 U3608 ( .A(n2147), .B(n4457), .Z(n3473) );
  AO4 U3609 ( .A(n3540), .B(n2666), .C(n3541), .D(n2577), .Z(n2271) );
  AO3 U3610 ( .A(n2264), .B(n2867), .C(n3542), .D(n3543), .Z(n3027) );
  AO2 U3611 ( .A(n2872), .B(n2268), .C(Datai[0]), .D(n2270), .Z(n3543) );
  IV U3612 ( .A(n2781), .Z(n2872) );
  ND2 U3613 ( .A(N2787), .B(n2364), .Z(n2781) );
  MUX21L U3614 ( .A(n2786), .B(n4409), .S(n2272), .Z(n3542) );
  AO4 U3615 ( .A(n3540), .B(n2645), .C(n3544), .D(n2577), .Z(n2786) );
  AO3 U3616 ( .A(n2264), .B(n2874), .C(n3545), .D(n3546), .Z(n3026) );
  AO2 U3617 ( .A(n2877), .B(n2268), .C(Datai[1]), .D(n2270), .Z(n3546) );
  IV U3618 ( .A(n2788), .Z(n2877) );
  ND2 U3619 ( .A(N2788), .B(n2364), .Z(n2788) );
  MUX21L U3620 ( .A(n2791), .B(n4421), .S(n2272), .Z(n3545) );
  AO4 U3621 ( .A(n3540), .B(n2648), .C(n3547), .D(n2577), .Z(n2791) );
  AO3 U3622 ( .A(n2264), .B(n2878), .C(n3548), .D(n3549), .Z(n3025) );
  AO2 U3623 ( .A(n2881), .B(n2268), .C(Datai[2]), .D(n2270), .Z(n3549) );
  IV U3624 ( .A(n2792), .Z(n2881) );
  ND2 U3625 ( .A(N2789), .B(n2364), .Z(n2792) );
  MUX21L U3626 ( .A(n2795), .B(n4399), .S(n2272), .Z(n3548) );
  AO4 U3627 ( .A(n3540), .B(n2651), .C(n3550), .D(n2577), .Z(n2795) );
  AO3 U3628 ( .A(n2264), .B(n2882), .C(n3551), .D(n3552), .Z(n3024) );
  AO2 U3629 ( .A(n2885), .B(n2268), .C(Datai[3]), .D(n2270), .Z(n3552) );
  IV U3630 ( .A(n2796), .Z(n2885) );
  ND2 U3631 ( .A(N2790), .B(n2364), .Z(n2796) );
  MUX21L U3632 ( .A(n2799), .B(n4432), .S(n2272), .Z(n3551) );
  AO4 U3633 ( .A(n3540), .B(n2654), .C(n3553), .D(n2577), .Z(n2799) );
  AO3 U3634 ( .A(n2264), .B(n2886), .C(n3554), .D(n3555), .Z(n3023) );
  AO2 U3635 ( .A(n2889), .B(n2268), .C(Datai[4]), .D(n2270), .Z(n3555) );
  IV U3636 ( .A(n2800), .Z(n2889) );
  ND2 U3637 ( .A(N2791), .B(n2364), .Z(n2800) );
  MUX21L U3638 ( .A(n2803), .B(n4442), .S(n2272), .Z(n3554) );
  AO4 U3639 ( .A(n3540), .B(n2657), .C(n3556), .D(n2577), .Z(n2803) );
  AO3 U3640 ( .A(n2264), .B(n2890), .C(n3557), .D(n3558), .Z(n3022) );
  AO2 U3641 ( .A(n2893), .B(n2268), .C(Datai[5]), .D(n2270), .Z(n3558) );
  IV U3642 ( .A(n2804), .Z(n2893) );
  ND2 U3643 ( .A(N2792), .B(n2364), .Z(n2804) );
  MUX21L U3644 ( .A(n2807), .B(n4368), .S(n2272), .Z(n3557) );
  AO4 U3645 ( .A(n3540), .B(n2660), .C(n3559), .D(n2577), .Z(n2807) );
  AO3 U3646 ( .A(n2264), .B(n2894), .C(n3560), .D(n3561), .Z(n3021) );
  AO2 U3647 ( .A(n2897), .B(n2268), .C(Datai[6]), .D(n2270), .Z(n3561) );
  NR4 U3648 ( .A(n2556), .B(n2272), .C(n2268), .D(n2816), .Z(n2270) );
  IV U3649 ( .A(n2808), .Z(n2897) );
  ND2 U3650 ( .A(N818), .B(n2364), .Z(n2808) );
  MUX21L U3651 ( .A(n2811), .B(n4389), .S(n2272), .Z(n3560) );
  NR3 U3652 ( .A(n2817), .B(n3538), .C(n3562), .Z(n2272) );
  AO4 U3653 ( .A(n2606), .B(n2820), .C(n2819), .D(n2822), .Z(n3562) );
  ND2 U3654 ( .A(n3332), .B(n3563), .Z(n2822) );
  NR2 U3655 ( .A(n2169), .B(n4455), .Z(n3332) );
  IV U3656 ( .A(n2276), .Z(n2819) );
  ND2 U3657 ( .A(n3356), .B(n3563), .Z(n2820) );
  NR2 U3658 ( .A(n4454), .B(n4455), .Z(n3356) );
  NR2 U3659 ( .A(n2276), .B(n2262), .Z(n2606) );
  IV U3660 ( .A(n2577), .Z(n2262) );
  IV U3661 ( .A(n3519), .Z(n3538) );
  ND2 U3662 ( .A(n2268), .B(n2364), .Z(n3519) );
  IV U3663 ( .A(n3496), .Z(n2268) );
  ND2 U3664 ( .A(n3563), .B(n3020), .Z(n3496) );
  NR2 U3665 ( .A(n2146), .B(n2169), .Z(n3020) );
  IV U3666 ( .A(n2264), .Z(n2817) );
  AO4 U3667 ( .A(n3540), .B(n2663), .C(n3564), .D(n2577), .Z(n2811) );
  ND3 U3668 ( .A(n2183), .B(n4668), .C(n3565), .Z(n2577) );
  ND2 U3669 ( .A(n2816), .B(n2364), .Z(n2264) );
  IV U3670 ( .A(n2780), .Z(n2816) );
  ND2 U3671 ( .A(n3308), .B(n3563), .Z(n2780) );
  NR2 U3672 ( .A(n4456), .B(n4457), .Z(n3563) );
  NR2 U3673 ( .A(n2146), .B(n4454), .Z(n3308) );
  AO7 U3674 ( .A(n4590), .B(n2626), .C(n3566), .Z(n3019) );
  AO2 U3675 ( .A(Datai[0]), .B(n2628), .C(N1750), .D(n2629), .Z(n3566) );
  AO7 U3676 ( .A(n4595), .B(n2626), .C(n3567), .Z(n3018) );
  AO2 U3677 ( .A(Datai[1]), .B(n2628), .C(N1751), .D(n2629), .Z(n3567) );
  AO7 U3678 ( .A(n4600), .B(n2626), .C(n3568), .Z(n3017) );
  AO2 U3679 ( .A(Datai[2]), .B(n2628), .C(N1752), .D(n2629), .Z(n3568) );
  AO7 U3680 ( .A(n4606), .B(n2626), .C(n3569), .Z(n3016) );
  AO2 U3681 ( .A(Datai[3]), .B(n2628), .C(N1753), .D(n2629), .Z(n3569) );
  AO7 U3682 ( .A(n4612), .B(n2626), .C(n3570), .Z(n3015) );
  AO2 U3683 ( .A(Datai[4]), .B(n2628), .C(N1754), .D(n2629), .Z(n3570) );
  AO7 U3684 ( .A(n4618), .B(n2626), .C(n3571), .Z(n3014) );
  AO2 U3685 ( .A(Datai[5]), .B(n2628), .C(N1755), .D(n2629), .Z(n3571) );
  AO7 U3686 ( .A(n4624), .B(n2626), .C(n3572), .Z(n3013) );
  AO2 U3687 ( .A(Datai[6]), .B(n2628), .C(N1756), .D(n2629), .Z(n3572) );
  AO7 U3688 ( .A(n4631), .B(n2626), .C(n3573), .Z(n3012) );
  AO2 U3689 ( .A(n2628), .B(Datai[7]), .C(n2629), .D(N1757), .Z(n3573) );
  AO7 U3690 ( .A(n4636), .B(n2626), .C(n3574), .Z(n3011) );
  AO2 U3691 ( .A(Datai[8]), .B(n2628), .C(N1758), .D(n2629), .Z(n3574) );
  AO7 U3692 ( .A(n4637), .B(n2626), .C(n3575), .Z(n3010) );
  AO2 U3693 ( .A(Datai[9]), .B(n2628), .C(N1759), .D(n2629), .Z(n3575) );
  AO7 U3694 ( .A(n4638), .B(n2626), .C(n3576), .Z(n3009) );
  AO2 U3695 ( .A(Datai[10]), .B(n2628), .C(N1760), .D(n2629), .Z(n3576) );
  AO7 U3696 ( .A(n4639), .B(n2626), .C(n3577), .Z(n3008) );
  AO2 U3697 ( .A(Datai[11]), .B(n2628), .C(N1761), .D(n2629), .Z(n3577) );
  AO7 U3698 ( .A(n4640), .B(n2626), .C(n3578), .Z(n3007) );
  AO2 U3699 ( .A(Datai[12]), .B(n2628), .C(N1762), .D(n2629), .Z(n3578) );
  AO7 U3700 ( .A(n4641), .B(n2626), .C(n3579), .Z(n3006) );
  AO2 U3701 ( .A(Datai[13]), .B(n2628), .C(N1763), .D(n2629), .Z(n3579) );
  AO7 U3702 ( .A(n4642), .B(n2626), .C(n3580), .Z(n3005) );
  AO2 U3703 ( .A(Datai[14]), .B(n2628), .C(N1764), .D(n2629), .Z(n3580) );
  NR2 U3704 ( .A(n2549), .B(n3581), .Z(n2629) );
  NR2 U3705 ( .A(n2395), .B(n3581), .Z(n2628) );
  IV U3706 ( .A(n2626), .Z(n3581) );
  AO7 U3707 ( .A(n2359), .B(n3582), .C(n3583), .Z(n2626) );
  MUX21L U3708 ( .A(n3584), .B(n4355), .S(n3585), .Z(n3004) );
  AO2 U3709 ( .A(n2371), .B(n2372), .C(n3586), .D(n3587), .Z(n3584) );
  AO3 U3710 ( .A(n2338), .B(n3588), .C(n3589), .D(n3590), .Z(n3003) );
  AO2 U3711 ( .A(n4654), .B(n2341), .C(rEIP[0]), .D(n2335), .Z(n3590) );
  ND2 U3712 ( .A(n317), .B(n2342), .Z(n3589) );
  IV U3713 ( .A(n460), .Z(n3588) );
  AO3 U3714 ( .A(n2338), .B(n3591), .C(n3592), .D(n3593), .Z(n3002) );
  AO2 U3715 ( .A(n4453), .B(n2341), .C(rEIP[1]), .D(n2335), .Z(n3593) );
  ND2 U3716 ( .A(n316), .B(n2342), .Z(n3592) );
  IV U3717 ( .A(n459), .Z(n3591) );
  AO3 U3718 ( .A(n2338), .B(n3594), .C(n3595), .D(n3596), .Z(n3001) );
  AO2 U3719 ( .A(n4473), .B(n2341), .C(rEIP[2]), .D(n2335), .Z(n3596) );
  ND2 U3720 ( .A(n315), .B(n2342), .Z(n3595) );
  IV U3721 ( .A(n458), .Z(n3594) );
  AO3 U3722 ( .A(n2338), .B(n3597), .C(n3598), .D(n3599), .Z(n3000) );
  AO2 U3723 ( .A(n4478), .B(n2341), .C(rEIP[3]), .D(n2335), .Z(n3599) );
  ND2 U3724 ( .A(n314), .B(n2342), .Z(n3598) );
  IV U3725 ( .A(n457), .Z(n3597) );
  AO3 U3726 ( .A(n2338), .B(n3600), .C(n3601), .D(n3602), .Z(n2999) );
  AO2 U3727 ( .A(n4483), .B(n2341), .C(rEIP[4]), .D(n2335), .Z(n3602) );
  ND2 U3728 ( .A(n313), .B(n2342), .Z(n3601) );
  IV U3729 ( .A(n456), .Z(n3600) );
  AO3 U3730 ( .A(n2338), .B(n3603), .C(n3604), .D(n3605), .Z(n2998) );
  AO2 U3731 ( .A(n4488), .B(n2341), .C(rEIP[5]), .D(n2335), .Z(n3605) );
  ND2 U3732 ( .A(n312), .B(n2342), .Z(n3604) );
  IV U3733 ( .A(n455), .Z(n3603) );
  AO3 U3734 ( .A(n2338), .B(n3606), .C(n3607), .D(n3608), .Z(n2997) );
  AO2 U3735 ( .A(n4493), .B(n2341), .C(rEIP[6]), .D(n2335), .Z(n3608) );
  ND2 U3736 ( .A(n311), .B(n2342), .Z(n3607) );
  IV U3737 ( .A(n454), .Z(n3606) );
  AO3 U3738 ( .A(n2338), .B(n3609), .C(n3610), .D(n3611), .Z(n2996) );
  AO2 U3739 ( .A(n4498), .B(n2341), .C(rEIP[7]), .D(n2335), .Z(n3611) );
  ND2 U3740 ( .A(n310), .B(n2342), .Z(n3610) );
  IV U3741 ( .A(n453), .Z(n3609) );
  AO3 U3742 ( .A(n2338), .B(n3612), .C(n3613), .D(n3614), .Z(n2995) );
  AO2 U3743 ( .A(n2341), .B(n2196), .C(rEIP[8]), .D(n2335), .Z(n3614) );
  ND2 U3744 ( .A(n309), .B(n2342), .Z(n3613) );
  IV U3745 ( .A(n452), .Z(n3612) );
  AO3 U3746 ( .A(n2338), .B(n3615), .C(n3616), .D(n3617), .Z(n2994) );
  AO2 U3747 ( .A(n2341), .B(n2195), .C(rEIP[9]), .D(n2335), .Z(n3617) );
  ND2 U3748 ( .A(n308), .B(n2342), .Z(n3616) );
  IV U3749 ( .A(n451), .Z(n3615) );
  AO3 U3750 ( .A(n2338), .B(n3618), .C(n3619), .D(n3620), .Z(n2993) );
  AO2 U3751 ( .A(n2341), .B(n2211), .C(rEIP[10]), .D(n2335), .Z(n3620) );
  ND2 U3752 ( .A(n307), .B(n2342), .Z(n3619) );
  IV U3753 ( .A(n450), .Z(n3618) );
  AO3 U3754 ( .A(n2338), .B(n3621), .C(n3622), .D(n3623), .Z(n2992) );
  AO2 U3755 ( .A(n2341), .B(n2210), .C(rEIP[11]), .D(n2335), .Z(n3623) );
  ND2 U3756 ( .A(n306), .B(n2342), .Z(n3622) );
  IV U3757 ( .A(n449), .Z(n3621) );
  AO3 U3758 ( .A(n2338), .B(n3624), .C(n3625), .D(n3626), .Z(n2991) );
  AO2 U3759 ( .A(n2341), .B(n2209), .C(rEIP[12]), .D(n2335), .Z(n3626) );
  ND2 U3760 ( .A(n305), .B(n2342), .Z(n3625) );
  IV U3761 ( .A(n448), .Z(n3624) );
  AO3 U3762 ( .A(n2338), .B(n3627), .C(n3628), .D(n3629), .Z(n2990) );
  AO2 U3763 ( .A(n2341), .B(n2208), .C(rEIP[13]), .D(n2335), .Z(n3629) );
  ND2 U3764 ( .A(n304), .B(n2342), .Z(n3628) );
  IV U3765 ( .A(n447), .Z(n3627) );
  AO3 U3766 ( .A(n2338), .B(n3630), .C(n3631), .D(n3632), .Z(n2989) );
  AO2 U3767 ( .A(n2341), .B(n2207), .C(rEIP[14]), .D(n2335), .Z(n3632) );
  ND2 U3768 ( .A(n303), .B(n2342), .Z(n3631) );
  IV U3769 ( .A(n446), .Z(n3630) );
  AO3 U3770 ( .A(n2338), .B(n3633), .C(n3634), .D(n3635), .Z(n2988) );
  AO2 U3771 ( .A(n2341), .B(n2206), .C(rEIP[15]), .D(n2335), .Z(n3635) );
  ND2 U3772 ( .A(n302), .B(n2342), .Z(n3634) );
  IV U3773 ( .A(n445), .Z(n3633) );
  AO3 U3774 ( .A(n2338), .B(n3636), .C(n3637), .D(n3638), .Z(n2987) );
  AO2 U3775 ( .A(n4536), .B(n2341), .C(rEIP[16]), .D(n2335), .Z(n3638) );
  ND2 U3776 ( .A(n301), .B(n2342), .Z(n3637) );
  AO3 U3777 ( .A(n2338), .B(n3639), .C(n3640), .D(n3641), .Z(n2986) );
  AO2 U3778 ( .A(n4540), .B(n2341), .C(rEIP[17]), .D(n2335), .Z(n3641) );
  ND2 U3779 ( .A(n300), .B(n2342), .Z(n3640) );
  AO3 U3780 ( .A(n2338), .B(n3642), .C(n3643), .D(n3644), .Z(n2985) );
  AO2 U3781 ( .A(n4544), .B(n2341), .C(rEIP[18]), .D(n2335), .Z(n3644) );
  ND2 U3782 ( .A(n299), .B(n2342), .Z(n3643) );
  AO3 U3783 ( .A(n2338), .B(n3645), .C(n3646), .D(n3647), .Z(n2984) );
  AO2 U3784 ( .A(n4548), .B(n2341), .C(rEIP[19]), .D(n2335), .Z(n3647) );
  ND2 U3785 ( .A(n298), .B(n2342), .Z(n3646) );
  IV U3786 ( .A(n441), .Z(n3645) );
  AO3 U3787 ( .A(n2338), .B(n3648), .C(n3649), .D(n3650), .Z(n2983) );
  AO2 U3788 ( .A(n4552), .B(n2341), .C(rEIP[20]), .D(n2335), .Z(n3650) );
  ND2 U3789 ( .A(n297), .B(n2342), .Z(n3649) );
  IV U3790 ( .A(n440), .Z(n3648) );
  AO3 U3791 ( .A(n2338), .B(n3651), .C(n3652), .D(n3653), .Z(n2982) );
  AO2 U3792 ( .A(n4556), .B(n2341), .C(rEIP[21]), .D(n2335), .Z(n3653) );
  ND2 U3793 ( .A(n296), .B(n2342), .Z(n3652) );
  IV U3794 ( .A(n439), .Z(n3651) );
  AO3 U3795 ( .A(n2338), .B(n3654), .C(n3655), .D(n3656), .Z(n2981) );
  AO2 U3796 ( .A(n4560), .B(n2341), .C(rEIP[22]), .D(n2335), .Z(n3656) );
  ND2 U3797 ( .A(n295), .B(n2342), .Z(n3655) );
  IV U3798 ( .A(n438), .Z(n3654) );
  AO3 U3799 ( .A(n2338), .B(n3657), .C(n3658), .D(n3659), .Z(n2980) );
  AO2 U3800 ( .A(n4564), .B(n2341), .C(rEIP[23]), .D(n2335), .Z(n3659) );
  ND2 U3801 ( .A(n294), .B(n2342), .Z(n3658) );
  AO3 U3802 ( .A(n2338), .B(n3660), .C(n3661), .D(n3662), .Z(n2979) );
  AO2 U3803 ( .A(n4568), .B(n2341), .C(rEIP[24]), .D(n2335), .Z(n3662) );
  ND2 U3804 ( .A(n293), .B(n2342), .Z(n3661) );
  AO3 U3805 ( .A(n2338), .B(n3663), .C(n3664), .D(n3665), .Z(n2978) );
  AO2 U3806 ( .A(n4572), .B(n2341), .C(rEIP[25]), .D(n2335), .Z(n3665) );
  ND2 U3807 ( .A(n292), .B(n2342), .Z(n3664) );
  AO3 U3808 ( .A(n2338), .B(n3666), .C(n3667), .D(n3668), .Z(n2977) );
  AO2 U3809 ( .A(n4576), .B(n2341), .C(rEIP[26]), .D(n2335), .Z(n3668) );
  ND2 U3810 ( .A(n291), .B(n2342), .Z(n3667) );
  AO3 U3811 ( .A(n2338), .B(n3669), .C(n3670), .D(n3671), .Z(n2976) );
  AO2 U3812 ( .A(n4580), .B(n2341), .C(rEIP[27]), .D(n2335), .Z(n3671) );
  ND2 U3813 ( .A(n290), .B(n2342), .Z(n3670) );
  AO3 U3814 ( .A(n2338), .B(n3672), .C(n3673), .D(n3674), .Z(n2975) );
  AO2 U3815 ( .A(n4584), .B(n2341), .C(rEIP[28]), .D(n2335), .Z(n3674) );
  ND2 U3816 ( .A(n289), .B(n2342), .Z(n3673) );
  AO3 U3817 ( .A(n2338), .B(n3675), .C(n3676), .D(n3677), .Z(n2974) );
  AO2 U3818 ( .A(n4588), .B(n2341), .C(rEIP[29]), .D(n2335), .Z(n3677) );
  ND2 U3819 ( .A(n288), .B(n2342), .Z(n3676) );
  AO3 U3820 ( .A(n2338), .B(n3678), .C(n3679), .D(n3680), .Z(n2973) );
  AO2 U3821 ( .A(n4645), .B(n2341), .C(rEIP[30]), .D(n2335), .Z(n3680) );
  ND2 U3822 ( .A(n287), .B(n2342), .Z(n3679) );
  NR3 U3823 ( .A(n2341), .B(n3681), .C(n2359), .Z(n2342) );
  NR4 U3824 ( .A(n2552), .B(n3682), .C(n3683), .D(n3684), .Z(n3681) );
  AO3 U3825 ( .A(n3685), .B(n3686), .C(n3687), .D(n2278), .Z(n2338) );
  IV U3826 ( .A(n2341), .Z(n3687) );
  NR3 U3827 ( .A(n2335), .B(n2580), .C(n3688), .Z(n2341) );
  NR2 U3828 ( .A(n2359), .B(n3689), .Z(n2580) );
  AN3 U3829 ( .A(n2616), .B(n3690), .C(n2615), .Z(n3689) );
  ND2 U3830 ( .A(n3691), .B(n2288), .Z(n2616) );
  ND2 U3831 ( .A(n2772), .B(n2549), .Z(n3686) );
  AO3 U3832 ( .A(n2332), .B(n3692), .C(n3693), .D(n3694), .Z(n2972) );
  AO2 U3833 ( .A(n460), .B(n2276), .C(rEIP[0]), .D(n2335), .Z(n3694) );
  OR2 U3834 ( .A(n2336), .B(n4460), .Z(n3693) );
  AO3 U3835 ( .A(n2332), .B(n3695), .C(n3696), .D(n3697), .Z(n2971) );
  AO2 U3836 ( .A(n459), .B(n2276), .C(rEIP[1]), .D(n2335), .Z(n3697) );
  OR2 U3837 ( .A(n2336), .B(n4459), .Z(n3696) );
  AO3 U3838 ( .A(n2332), .B(n3698), .C(n3699), .D(n3700), .Z(n2970) );
  AO2 U3839 ( .A(n458), .B(n2276), .C(rEIP[2]), .D(n2335), .Z(n3700) );
  OR2 U3840 ( .A(n2336), .B(n4472), .Z(n3699) );
  AO3 U3841 ( .A(n2332), .B(n3701), .C(n3702), .D(n3703), .Z(n2969) );
  AO2 U3842 ( .A(n457), .B(n2276), .C(rEIP[3]), .D(n2335), .Z(n3703) );
  OR2 U3843 ( .A(n2336), .B(n4477), .Z(n3702) );
  AO3 U3844 ( .A(n2332), .B(n3704), .C(n3705), .D(n3706), .Z(n2968) );
  AO2 U3845 ( .A(n456), .B(n2276), .C(rEIP[4]), .D(n2335), .Z(n3706) );
  ND2 U3846 ( .A(n2370), .B(n2185), .Z(n3705) );
  AO3 U3847 ( .A(n2332), .B(n3707), .C(n3708), .D(n3709), .Z(n2967) );
  AO2 U3848 ( .A(n455), .B(n2276), .C(rEIP[5]), .D(n2335), .Z(n3709) );
  ND2 U3849 ( .A(n2370), .B(n2186), .Z(n3708) );
  IV U3850 ( .A(n2336), .Z(n2370) );
  AO3 U3851 ( .A(n2332), .B(n2436), .C(n3710), .D(n3711), .Z(n2966) );
  AO2 U3852 ( .A(n454), .B(n2276), .C(rEIP[6]), .D(n2335), .Z(n3711) );
  OR2 U3853 ( .A(n2336), .B(n4492), .Z(n3710) );
  AO3 U3854 ( .A(n2332), .B(n2441), .C(n3712), .D(n3713), .Z(n2965) );
  AO2 U3855 ( .A(n453), .B(n2276), .C(rEIP[7]), .D(n2335), .Z(n3713) );
  OR2 U3856 ( .A(n2336), .B(n4497), .Z(n3712) );
  AO3 U3857 ( .A(n2332), .B(n2446), .C(n3714), .D(n3715), .Z(n2964) );
  AO2 U3858 ( .A(n452), .B(n2276), .C(rEIP[8]), .D(n2335), .Z(n3715) );
  OR2 U3859 ( .A(n2336), .B(n4502), .Z(n3714) );
  AO3 U3860 ( .A(n2332), .B(n2451), .C(n3716), .D(n3717), .Z(n2963) );
  AO2 U3861 ( .A(n451), .B(n2276), .C(rEIP[9]), .D(n2335), .Z(n3717) );
  OR2 U3862 ( .A(n2336), .B(n4506), .Z(n3716) );
  AO3 U3863 ( .A(n2332), .B(n2456), .C(n3718), .D(n3719), .Z(n2962) );
  AO2 U3864 ( .A(n450), .B(n2276), .C(rEIP[10]), .D(n2335), .Z(n3719) );
  OR2 U3865 ( .A(n2336), .B(n4510), .Z(n3718) );
  AO3 U3866 ( .A(n2332), .B(n2461), .C(n3720), .D(n3721), .Z(n2961) );
  AO2 U3867 ( .A(n449), .B(n2276), .C(rEIP[11]), .D(n2335), .Z(n3721) );
  OR2 U3868 ( .A(n2336), .B(n4514), .Z(n3720) );
  AO3 U3869 ( .A(n2332), .B(n2466), .C(n3722), .D(n3723), .Z(n2960) );
  AO2 U3870 ( .A(n448), .B(n2276), .C(rEIP[12]), .D(n2335), .Z(n3723) );
  OR2 U3871 ( .A(n2336), .B(n4518), .Z(n3722) );
  AO3 U3872 ( .A(n2332), .B(n2471), .C(n3724), .D(n3725), .Z(n2959) );
  AO2 U3873 ( .A(n447), .B(n2276), .C(rEIP[13]), .D(n2335), .Z(n3725) );
  OR2 U3874 ( .A(n2336), .B(n4522), .Z(n3724) );
  AO3 U3875 ( .A(n2332), .B(n2476), .C(n3726), .D(n3727), .Z(n2958) );
  AO2 U3876 ( .A(n446), .B(n2276), .C(rEIP[14]), .D(n2335), .Z(n3727) );
  OR2 U3877 ( .A(n2336), .B(n4526), .Z(n3726) );
  AO3 U3878 ( .A(n2332), .B(n2481), .C(n3728), .D(n3729), .Z(n2957) );
  AO2 U3879 ( .A(n445), .B(n2276), .C(rEIP[15]), .D(n2335), .Z(n3729) );
  OR2 U3880 ( .A(n2336), .B(n4530), .Z(n3728) );
  AO3 U3881 ( .A(n2332), .B(n2486), .C(n3730), .D(n3731), .Z(n2956) );
  AO2 U3882 ( .A(n444), .B(n2276), .C(rEIP[16]), .D(n2335), .Z(n3731) );
  OR2 U3883 ( .A(n2336), .B(n4535), .Z(n3730) );
  AO3 U3884 ( .A(n2332), .B(n2491), .C(n3732), .D(n3733), .Z(n2955) );
  AO2 U3885 ( .A(n443), .B(n2276), .C(rEIP[17]), .D(n2335), .Z(n3733) );
  OR2 U3886 ( .A(n2336), .B(n4539), .Z(n3732) );
  AO3 U3887 ( .A(n2332), .B(n2496), .C(n3734), .D(n3735), .Z(n2954) );
  AO2 U3888 ( .A(n442), .B(n2276), .C(rEIP[18]), .D(n2335), .Z(n3735) );
  OR2 U3889 ( .A(n2336), .B(n4543), .Z(n3734) );
  AO3 U3890 ( .A(n2332), .B(n2501), .C(n3736), .D(n3737), .Z(n2953) );
  AO2 U3891 ( .A(n441), .B(n2276), .C(rEIP[19]), .D(n2335), .Z(n3737) );
  OR2 U3892 ( .A(n2336), .B(n4547), .Z(n3736) );
  AO3 U3893 ( .A(n2332), .B(n2505), .C(n3738), .D(n3739), .Z(n2952) );
  AO2 U3894 ( .A(n440), .B(n2276), .C(rEIP[20]), .D(n2335), .Z(n3739) );
  OR2 U3895 ( .A(n2336), .B(n4551), .Z(n3738) );
  AO3 U3896 ( .A(n2332), .B(n2509), .C(n3740), .D(n3741), .Z(n2951) );
  AO2 U3897 ( .A(n439), .B(n2276), .C(rEIP[21]), .D(n2335), .Z(n3741) );
  OR2 U3898 ( .A(n2336), .B(n4555), .Z(n3740) );
  AO3 U3899 ( .A(n2332), .B(n2513), .C(n3742), .D(n3743), .Z(n2950) );
  AO2 U3900 ( .A(n438), .B(n2276), .C(rEIP[22]), .D(n2335), .Z(n3743) );
  OR2 U3901 ( .A(n2336), .B(n4559), .Z(n3742) );
  AO3 U3902 ( .A(n2332), .B(n2517), .C(n3744), .D(n3745), .Z(n2949) );
  AO2 U3903 ( .A(n437), .B(n2276), .C(rEIP[23]), .D(n2335), .Z(n3745) );
  OR2 U3904 ( .A(n2336), .B(n4563), .Z(n3744) );
  AO3 U3905 ( .A(n2332), .B(n2521), .C(n3746), .D(n3747), .Z(n2948) );
  AO2 U3906 ( .A(n436), .B(n2276), .C(rEIP[24]), .D(n2335), .Z(n3747) );
  OR2 U3907 ( .A(n2336), .B(n4567), .Z(n3746) );
  AO3 U3908 ( .A(n2332), .B(n2525), .C(n3748), .D(n3749), .Z(n2947) );
  AO2 U3909 ( .A(n435), .B(n2276), .C(rEIP[25]), .D(n2335), .Z(n3749) );
  OR2 U3910 ( .A(n2336), .B(n4571), .Z(n3748) );
  AO3 U3911 ( .A(n2332), .B(n2529), .C(n3750), .D(n3751), .Z(n2946) );
  AO2 U3912 ( .A(n434), .B(n2276), .C(rEIP[26]), .D(n2335), .Z(n3751) );
  OR2 U3913 ( .A(n2336), .B(n4575), .Z(n3750) );
  AO3 U3914 ( .A(n2332), .B(n2533), .C(n3752), .D(n3753), .Z(n2945) );
  AO2 U3915 ( .A(n433), .B(n2276), .C(rEIP[27]), .D(n2335), .Z(n3753) );
  OR2 U3916 ( .A(n2336), .B(n4579), .Z(n3752) );
  AO3 U3917 ( .A(n2332), .B(n2537), .C(n3754), .D(n3755), .Z(n2944) );
  AO2 U3918 ( .A(n432), .B(n2276), .C(rEIP[28]), .D(n2335), .Z(n3755) );
  OR2 U3919 ( .A(n2336), .B(n4583), .Z(n3754) );
  AO3 U3920 ( .A(n2332), .B(n2541), .C(n3756), .D(n3757), .Z(n2943) );
  AO2 U3921 ( .A(n431), .B(n2276), .C(rEIP[29]), .D(n2335), .Z(n3757) );
  OR2 U3922 ( .A(n2336), .B(n4587), .Z(n3756) );
  AO3 U3923 ( .A(n2332), .B(n2545), .C(n3758), .D(n3759), .Z(n2942) );
  AO2 U3924 ( .A(n430), .B(n2276), .C(rEIP[30]), .D(n2335), .Z(n3759) );
  OR2 U3925 ( .A(n2336), .B(n4644), .Z(n3758) );
  ND2 U3926 ( .A(n2278), .B(n2336), .Z(n2332) );
  OR3 U3927 ( .A(n3688), .B(n2335), .C(n2276), .Z(n2336) );
  ND2 U3928 ( .A(n2556), .B(n2360), .Z(n2276) );
  NR2 U3929 ( .A(n3760), .B(n2396), .Z(n2335) );
  NR2 U3930 ( .A(n2359), .B(n3761), .Z(n3688) );
  AO7 U3931 ( .A(n5315), .B(n3762), .C(n3763), .Z(n2941) );
  AO2 U3932 ( .A(n3764), .B(n4465), .C(n3765), .D(n234), .Z(n3763) );
  AO7 U3933 ( .A(n5314), .B(n3762), .C(n3766), .Z(n2940) );
  AO2 U3934 ( .A(n3764), .B(n4469), .C(n3765), .D(n233), .Z(n3766) );
  AO7 U3935 ( .A(n5313), .B(n3762), .C(n3767), .Z(n2939) );
  AO2 U3936 ( .A(n3764), .B(n4474), .C(n3765), .D(n232), .Z(n3767) );
  AO7 U3937 ( .A(n5312), .B(n3762), .C(n3768), .Z(n2938) );
  AO2 U3938 ( .A(n3764), .B(n4479), .C(n3765), .D(n231), .Z(n3768) );
  AO7 U3939 ( .A(n5311), .B(n3762), .C(n3769), .Z(n2937) );
  AO2 U3940 ( .A(n3764), .B(n4484), .C(n3765), .D(n230), .Z(n3769) );
  AO7 U3941 ( .A(n5310), .B(n3762), .C(n3770), .Z(n2936) );
  AO2 U3942 ( .A(n3764), .B(n4489), .C(n3765), .D(n229), .Z(n3770) );
  AO7 U3943 ( .A(n5309), .B(n3762), .C(n3771), .Z(n2935) );
  AO2 U3944 ( .A(n3764), .B(n4494), .C(n3765), .D(n228), .Z(n3771) );
  AO7 U3945 ( .A(n5308), .B(n3762), .C(n3772), .Z(n2934) );
  AO2 U3946 ( .A(n3764), .B(n4499), .C(n3765), .D(n227), .Z(n3772) );
  AO7 U3947 ( .A(n5307), .B(n3762), .C(n3773), .Z(n2933) );
  AO2 U3948 ( .A(n3764), .B(n4503), .C(n3765), .D(n226), .Z(n3773) );
  AO7 U3949 ( .A(n5306), .B(n3762), .C(n3774), .Z(n2932) );
  AO2 U3950 ( .A(n3764), .B(n4507), .C(n3765), .D(n225), .Z(n3774) );
  AO7 U3951 ( .A(n5305), .B(n3762), .C(n3775), .Z(n2931) );
  AO2 U3952 ( .A(n3764), .B(n4511), .C(n3765), .D(n224), .Z(n3775) );
  AO7 U3953 ( .A(n5304), .B(n3762), .C(n3776), .Z(n2930) );
  AO2 U3954 ( .A(n3764), .B(n4515), .C(n3765), .D(n223), .Z(n3776) );
  AO7 U3955 ( .A(n5303), .B(n3762), .C(n3777), .Z(n2929) );
  AO2 U3956 ( .A(n3764), .B(n4519), .C(n3765), .D(n222), .Z(n3777) );
  AO7 U3957 ( .A(n5302), .B(n3762), .C(n3778), .Z(n2928) );
  AO2 U3958 ( .A(n3764), .B(n4523), .C(n3765), .D(n221), .Z(n3778) );
  AO7 U3959 ( .A(n5301), .B(n3762), .C(n3779), .Z(n2927) );
  AO2 U3960 ( .A(n3764), .B(n4527), .C(n3765), .D(n220), .Z(n3779) );
  AO7 U3961 ( .A(n5300), .B(n3762), .C(n3780), .Z(n2926) );
  AO2 U3962 ( .A(n3764), .B(n4531), .C(n3765), .D(n219), .Z(n3780) );
  NR3 U3963 ( .A(n2359), .B(n3781), .C(n2283), .Z(n3764) );
  AO4 U3964 ( .A(n5426), .B(n3762), .C(n2485), .D(n3782), .Z(n2925) );
  AO4 U3965 ( .A(n5425), .B(n3762), .C(n2490), .D(n3782), .Z(n2924) );
  AO4 U3966 ( .A(n5424), .B(n3762), .C(n2495), .D(n3782), .Z(n2923) );
  AO4 U3967 ( .A(n5423), .B(n3762), .C(n2500), .D(n3782), .Z(n2922) );
  AO4 U3968 ( .A(n5422), .B(n3762), .C(n3783), .D(n3782), .Z(n2921) );
  AO4 U3969 ( .A(n5421), .B(n3762), .C(n3784), .D(n3782), .Z(n2920) );
  AO4 U3970 ( .A(n5420), .B(n3762), .C(n3785), .D(n3782), .Z(n2919) );
  AO4 U3971 ( .A(n5419), .B(n3762), .C(n3786), .D(n3782), .Z(n2918) );
  AO4 U3972 ( .A(n5418), .B(n3762), .C(n3787), .D(n3782), .Z(n2917) );
  AO4 U3973 ( .A(n5417), .B(n3762), .C(n3788), .D(n3782), .Z(n2916) );
  AO4 U3974 ( .A(n5416), .B(n3762), .C(n3789), .D(n3782), .Z(n2915) );
  AO4 U3975 ( .A(n5415), .B(n3762), .C(n3790), .D(n3782), .Z(n2914) );
  AO4 U3976 ( .A(n5414), .B(n3762), .C(n3791), .D(n3782), .Z(n2913) );
  AO4 U3977 ( .A(n5413), .B(n3762), .C(n3792), .D(n3782), .Z(n2912) );
  AO4 U3978 ( .A(n5412), .B(n3762), .C(n3793), .D(n3782), .Z(n2911) );
  IV U3979 ( .A(n3765), .Z(n3782) );
  AO6 U3980 ( .A(n2549), .B(n2357), .C(n3781), .Z(n3765) );
  IV U3981 ( .A(n3762), .Z(n3781) );
  AO3 U3982 ( .A(n2283), .B(n3794), .C(n2357), .D(n3795), .Z(n3762) );
  ND2 U3983 ( .A(n3796), .B(n2284), .Z(n3794) );
  AO3 U3984 ( .A(n4648), .B(n3797), .C(n3798), .D(n3799), .Z(n2910) );
  ND2 U3985 ( .A(n4656), .B(n2149), .Z(n3799) );
  MUX21L U3986 ( .A(n5411), .B(n4648), .S(n2246), .Z(n2909) );
  AO3 U3987 ( .A(n2168), .B(n3800), .C(n3801), .D(n3802), .Z(n2908) );
  OR2 U3988 ( .A(n3797), .B(n4356), .Z(n3802) );
  AO3 U3989 ( .A(n4655), .B(n2168), .C(n2149), .D(n4656), .Z(n3801) );
  AO3 U3990 ( .A(n4649), .B(n3797), .C(n3800), .D(n3798), .Z(n2907) );
  ND3 U3991 ( .A(n2168), .B(n4656), .C(n4655), .Z(n3798) );
  ND2 U3992 ( .A(n3803), .B(n3800), .Z(n2906) );
  ND2 U3993 ( .A(rEIP[1]), .B(n3797), .Z(n3800) );
  MUX21H U3994 ( .A(n4650), .B(n2168), .S(n3797), .Z(n3803) );
  OR2 U3995 ( .A(n4655), .B(n4656), .Z(n3797) );
  MUX21L U3996 ( .A(n5409), .B(n4650), .S(n2246), .Z(n2905) );
  MUX21L U3997 ( .A(n3761), .B(n4357), .S(n3585), .Z(n22) );
  ND2 U3998 ( .A(n2278), .B(n2386), .Z(n3585) );
  ND4 U3999 ( .A(n3804), .B(n3805), .C(n3806), .D(n2387), .Z(n2386) );
  ND2 U4000 ( .A(n2286), .B(n3807), .Z(n3806) );
  ND3 U4001 ( .A(n3808), .B(n2395), .C(n2287), .Z(n3807) );
  NR2 U4002 ( .A(n3809), .B(n3810), .Z(n3761) );
  AO3 U4003 ( .A(n3811), .B(n3812), .C(n3813), .D(n3814), .Z(n2144) );
  AO2 U4004 ( .A(n3815), .B(n441), .C(n3816), .D(n3817), .Z(n3814) );
  ND2 U4005 ( .A(n3818), .B(n2187), .Z(n3813) );
  AO6 U4006 ( .A(n3819), .B(n3820), .C(n3821), .Z(n3811) );
  AO4 U4007 ( .A(n2570), .B(n3822), .C(n4468), .D(n3823), .Z(n3821) );
  AO7 U4008 ( .A(n3642), .B(n3824), .C(n3825), .Z(n2143) );
  AO2 U4009 ( .A(n3826), .B(n3827), .C(n3818), .D(n2188), .Z(n3825) );
  AO7 U4010 ( .A(n2610), .B(n3828), .C(n3829), .Z(n3827) );
  EO1 U4011 ( .A(n3830), .B(n2145), .C(n3831), .D(n2570), .Z(n3829) );
  IV U4012 ( .A(n442), .Z(n3642) );
  AO7 U4013 ( .A(n3639), .B(n3824), .C(n3832), .Z(n2142) );
  AO2 U4014 ( .A(n3826), .B(n3833), .C(n3818), .D(n2189), .Z(n3832) );
  AO7 U4015 ( .A(n2610), .B(n3834), .C(n3835), .Z(n3833) );
  EO1 U4016 ( .A(n3836), .B(n2145), .C(n3837), .D(n2570), .Z(n3835) );
  IV U4017 ( .A(n443), .Z(n3639) );
  AO7 U4018 ( .A(n3636), .B(n3824), .C(n3838), .Z(n2141) );
  AO2 U4019 ( .A(n3826), .B(n3839), .C(n3818), .D(n2190), .Z(n3838) );
  IV U4020 ( .A(n3840), .Z(n3818) );
  AO7 U4021 ( .A(n2610), .B(n3841), .C(n3842), .Z(n3839) );
  AO2 U4022 ( .A(n3843), .B(n2145), .C(n3844), .D(n2573), .Z(n3842) );
  IV U4023 ( .A(n444), .Z(n3636) );
  AO7 U4024 ( .A(n2590), .B(n2751), .C(n3845), .Z(n2140) );
  IV U4025 ( .A(Datai[24]), .Z(n2751) );
  NR2 U4026 ( .A(n2590), .B(n2775), .Z(U3_U8_Z_7) );
  NR2 U4027 ( .A(n2590), .B(n2769), .Z(U3_U8_Z_6) );
  IV U4028 ( .A(Datai[30]), .Z(n2769) );
  NR2 U4029 ( .A(n2590), .B(n2766), .Z(U3_U8_Z_5) );
  IV U4030 ( .A(Datai[29]), .Z(n2766) );
  NR2 U4031 ( .A(n2590), .B(n2763), .Z(U3_U8_Z_4) );
  IV U4032 ( .A(Datai[28]), .Z(n2763) );
  NR2 U4033 ( .A(n2590), .B(n2760), .Z(U3_U8_Z_3) );
  IV U4034 ( .A(Datai[27]), .Z(n2760) );
  NR2 U4035 ( .A(n2590), .B(n2757), .Z(U3_U8_Z_2) );
  IV U4036 ( .A(Datai[26]), .Z(n2757) );
  NR2 U4037 ( .A(n2590), .B(n2754), .Z(U3_U8_Z_1) );
  IV U4038 ( .A(Datai[25]), .Z(n2754) );
  NR2 U4039 ( .A(n4467), .B(n3845), .Z(U3_U7_Z_3) );
  NR2 U4040 ( .A(n4653), .B(n3845), .Z(U3_U7_Z_2) );
  NR2 U4041 ( .A(n4461), .B(n3845), .Z(U3_U7_Z_1) );
  AO4 U4042 ( .A(n4468), .B(n3845), .C(n3846), .D(n2590), .Z(U3_U7_Z_0) );
  NR2 U4043 ( .A(n3847), .B(n3848), .Z(n3846) );
  AO6 U4044 ( .A(n3849), .B(n3850), .C(n2775), .Z(n3848) );
  IV U4045 ( .A(Datai[31]), .Z(n2775) );
  NR4 U4046 ( .A(Datai[23]), .B(Datai[22]), .C(Datai[21]), .D(Datai[20]), .Z(
        n3850) );
  NR4 U4047 ( .A(Datai[19]), .B(Datai[18]), .C(Datai[17]), .D(Datai[16]), .Z(
        n3849) );
  IV U4048 ( .A(n3851), .Z(n3847) );
  ND2 U4049 ( .A(n3796), .B(n3684), .Z(n3845) );
  AO4 U4050 ( .A(n2615), .B(n2451), .C(n3582), .D(n2672), .Z(U3_U6_Z_9) );
  IV U4051 ( .A(n308), .Z(n2451) );
  AO4 U4052 ( .A(n2615), .B(n2446), .C(n3582), .D(n2669), .Z(U3_U6_Z_8) );
  IV U4053 ( .A(n309), .Z(n2446) );
  AO4 U4054 ( .A(n2615), .B(n2441), .C(n2666), .D(n3582), .Z(U3_U6_Z_7) );
  IV U4055 ( .A(n310), .Z(n2441) );
  AO4 U4056 ( .A(n2615), .B(n2436), .C(n3582), .D(n2663), .Z(U3_U6_Z_6) );
  IV U4057 ( .A(n311), .Z(n2436) );
  AO4 U4058 ( .A(n2615), .B(n3707), .C(n3582), .D(n2660), .Z(U3_U6_Z_5) );
  IV U4059 ( .A(n312), .Z(n3707) );
  AO4 U4060 ( .A(n2615), .B(n3704), .C(n3582), .D(n2657), .Z(U3_U6_Z_4) );
  IV U4061 ( .A(n313), .Z(n3704) );
  NR2 U4062 ( .A(n2615), .B(n2545), .Z(U3_U6_Z_30) );
  IV U4063 ( .A(n287), .Z(n2545) );
  AO4 U4064 ( .A(n2615), .B(n3701), .C(n3582), .D(n2654), .Z(U3_U6_Z_3) );
  IV U4065 ( .A(n314), .Z(n3701) );
  NR2 U4066 ( .A(n2615), .B(n2541), .Z(U3_U6_Z_29) );
  IV U4067 ( .A(n288), .Z(n2541) );
  NR2 U4068 ( .A(n2615), .B(n2537), .Z(U3_U6_Z_28) );
  IV U4069 ( .A(n289), .Z(n2537) );
  NR2 U4070 ( .A(n2615), .B(n2533), .Z(U3_U6_Z_27) );
  IV U4071 ( .A(n290), .Z(n2533) );
  NR2 U4072 ( .A(n2615), .B(n2529), .Z(U3_U6_Z_26) );
  IV U4073 ( .A(n291), .Z(n2529) );
  NR2 U4074 ( .A(n2615), .B(n2525), .Z(U3_U6_Z_25) );
  IV U4075 ( .A(n292), .Z(n2525) );
  NR2 U4076 ( .A(n2615), .B(n2521), .Z(U3_U6_Z_24) );
  IV U4077 ( .A(n293), .Z(n2521) );
  NR2 U4078 ( .A(n2615), .B(n2517), .Z(U3_U6_Z_23) );
  IV U4079 ( .A(n294), .Z(n2517) );
  NR2 U4080 ( .A(n2615), .B(n2513), .Z(U3_U6_Z_22) );
  IV U4081 ( .A(n295), .Z(n2513) );
  NR2 U4082 ( .A(n2615), .B(n2509), .Z(U3_U6_Z_21) );
  IV U4083 ( .A(n296), .Z(n2509) );
  NR2 U4084 ( .A(n2615), .B(n2505), .Z(U3_U6_Z_20) );
  IV U4085 ( .A(n297), .Z(n2505) );
  AO4 U4086 ( .A(n2615), .B(n3698), .C(n3582), .D(n2651), .Z(U3_U6_Z_2) );
  IV U4087 ( .A(n315), .Z(n3698) );
  NR2 U4088 ( .A(n2615), .B(n2501), .Z(U3_U6_Z_19) );
  IV U4089 ( .A(n298), .Z(n2501) );
  NR2 U4090 ( .A(n2615), .B(n2496), .Z(U3_U6_Z_18) );
  IV U4091 ( .A(n299), .Z(n2496) );
  NR2 U4092 ( .A(n2615), .B(n2491), .Z(U3_U6_Z_17) );
  IV U4093 ( .A(n300), .Z(n2491) );
  NR2 U4094 ( .A(n2615), .B(n2486), .Z(U3_U6_Z_16) );
  IV U4095 ( .A(n301), .Z(n2486) );
  AO4 U4096 ( .A(n2615), .B(n2481), .C(n2620), .D(n3582), .Z(U3_U6_Z_15) );
  IV U4097 ( .A(Datai[15]), .Z(n2620) );
  IV U4098 ( .A(n302), .Z(n2481) );
  AO4 U4099 ( .A(n2615), .B(n2476), .C(n3582), .D(n2687), .Z(U3_U6_Z_14) );
  IV U4100 ( .A(n303), .Z(n2476) );
  AO4 U4101 ( .A(n2615), .B(n2471), .C(n3582), .D(n2684), .Z(U3_U6_Z_13) );
  IV U4102 ( .A(n304), .Z(n2471) );
  AO4 U4103 ( .A(n2615), .B(n2466), .C(n3582), .D(n2681), .Z(U3_U6_Z_12) );
  IV U4104 ( .A(n305), .Z(n2466) );
  AO4 U4105 ( .A(n2615), .B(n2461), .C(n3582), .D(n2678), .Z(U3_U6_Z_11) );
  IV U4106 ( .A(n306), .Z(n2461) );
  AO4 U4107 ( .A(n2615), .B(n2456), .C(n3582), .D(n2675), .Z(U3_U6_Z_10) );
  IV U4108 ( .A(n307), .Z(n2456) );
  AO4 U4109 ( .A(n2615), .B(n3695), .C(n3582), .D(n2648), .Z(U3_U6_Z_1) );
  IV U4110 ( .A(n316), .Z(n3695) );
  AO4 U4111 ( .A(n2615), .B(n3692), .C(n3582), .D(n2645), .Z(U3_U6_Z_0) );
  IV U4112 ( .A(n317), .Z(n3692) );
  NR2 U4113 ( .A(n2615), .B(n2450), .Z(U3_U5_Z_9) );
  IV U4114 ( .A(n225), .Z(n2450) );
  NR2 U4115 ( .A(n2615), .B(n2445), .Z(U3_U5_Z_8) );
  IV U4116 ( .A(n226), .Z(n2445) );
  NR2 U4117 ( .A(n2615), .B(n2440), .Z(U3_U5_Z_7) );
  IV U4118 ( .A(n227), .Z(n2440) );
  NR2 U4119 ( .A(n2615), .B(n2435), .Z(U3_U5_Z_6) );
  IV U4120 ( .A(n228), .Z(n2435) );
  AN2 U4121 ( .A(n2613), .B(n229), .Z(U3_U5_Z_5) );
  AN2 U4122 ( .A(n2613), .B(n230), .Z(U3_U5_Z_4) );
  AO4 U4123 ( .A(n2615), .B(n3793), .C(n3582), .D(n2687), .Z(U3_U5_Z_30) );
  IV U4124 ( .A(Datai[14]), .Z(n2687) );
  IV U4125 ( .A(n204), .Z(n3793) );
  AN2 U4126 ( .A(n2613), .B(n231), .Z(U3_U5_Z_3) );
  AO4 U4127 ( .A(n2615), .B(n3792), .C(n3582), .D(n2684), .Z(U3_U5_Z_29) );
  IV U4128 ( .A(Datai[13]), .Z(n2684) );
  IV U4129 ( .A(n205), .Z(n3792) );
  AO4 U4130 ( .A(n2615), .B(n3791), .C(n3582), .D(n2681), .Z(U3_U5_Z_28) );
  IV U4131 ( .A(Datai[12]), .Z(n2681) );
  IV U4132 ( .A(n206), .Z(n3791) );
  AO4 U4133 ( .A(n2615), .B(n3790), .C(n3582), .D(n2678), .Z(U3_U5_Z_27) );
  IV U4134 ( .A(Datai[11]), .Z(n2678) );
  IV U4135 ( .A(n207), .Z(n3790) );
  AO4 U4136 ( .A(n2615), .B(n3789), .C(n3582), .D(n2675), .Z(U3_U5_Z_26) );
  IV U4137 ( .A(Datai[10]), .Z(n2675) );
  IV U4138 ( .A(n208), .Z(n3789) );
  AO4 U4139 ( .A(n2615), .B(n3788), .C(n3582), .D(n2672), .Z(U3_U5_Z_25) );
  IV U4140 ( .A(Datai[9]), .Z(n2672) );
  IV U4141 ( .A(n209), .Z(n3788) );
  AO4 U4142 ( .A(n2615), .B(n3787), .C(n3582), .D(n2669), .Z(U3_U5_Z_24) );
  IV U4143 ( .A(Datai[8]), .Z(n2669) );
  IV U4144 ( .A(n210), .Z(n3787) );
  AO4 U4145 ( .A(n2615), .B(n3786), .C(n2666), .D(n3582), .Z(U3_U5_Z_23) );
  IV U4146 ( .A(Datai[7]), .Z(n2666) );
  IV U4147 ( .A(n211), .Z(n3786) );
  AO4 U4148 ( .A(n2615), .B(n3785), .C(n3582), .D(n2663), .Z(U3_U5_Z_22) );
  IV U4149 ( .A(Datai[6]), .Z(n2663) );
  IV U4150 ( .A(n212), .Z(n3785) );
  AO4 U4151 ( .A(n2615), .B(n3784), .C(n3582), .D(n2660), .Z(U3_U5_Z_21) );
  IV U4152 ( .A(Datai[5]), .Z(n2660) );
  IV U4153 ( .A(n213), .Z(n3784) );
  AO4 U4154 ( .A(n2615), .B(n3783), .C(n3582), .D(n2657), .Z(U3_U5_Z_20) );
  IV U4155 ( .A(Datai[4]), .Z(n2657) );
  IV U4156 ( .A(n214), .Z(n3783) );
  AN2 U4157 ( .A(n2613), .B(n232), .Z(U3_U5_Z_2) );
  AO4 U4158 ( .A(n2615), .B(n2500), .C(n3582), .D(n2654), .Z(U3_U5_Z_19) );
  IV U4159 ( .A(Datai[3]), .Z(n2654) );
  IV U4160 ( .A(n215), .Z(n2500) );
  AO4 U4161 ( .A(n2615), .B(n2495), .C(n3582), .D(n2651), .Z(U3_U5_Z_18) );
  IV U4162 ( .A(Datai[2]), .Z(n2651) );
  IV U4163 ( .A(n216), .Z(n2495) );
  AO4 U4164 ( .A(n2615), .B(n2490), .C(n3582), .D(n2648), .Z(U3_U5_Z_17) );
  IV U4165 ( .A(Datai[1]), .Z(n2648) );
  IV U4166 ( .A(n217), .Z(n2490) );
  AO4 U4167 ( .A(n2615), .B(n2485), .C(n3582), .D(n2645), .Z(U3_U5_Z_16) );
  IV U4168 ( .A(Datai[0]), .Z(n2645) );
  IV U4169 ( .A(n218), .Z(n2485) );
  NR2 U4170 ( .A(n2615), .B(n2480), .Z(U3_U5_Z_15) );
  IV U4171 ( .A(n219), .Z(n2480) );
  NR2 U4172 ( .A(n2615), .B(n2475), .Z(U3_U5_Z_14) );
  IV U4173 ( .A(n220), .Z(n2475) );
  NR2 U4174 ( .A(n2615), .B(n2470), .Z(U3_U5_Z_13) );
  IV U4175 ( .A(n221), .Z(n2470) );
  NR2 U4176 ( .A(n2615), .B(n2465), .Z(U3_U5_Z_12) );
  IV U4177 ( .A(n222), .Z(n2465) );
  NR2 U4178 ( .A(n2615), .B(n2460), .Z(U3_U5_Z_11) );
  IV U4179 ( .A(n223), .Z(n2460) );
  NR2 U4180 ( .A(n2615), .B(n2455), .Z(U3_U5_Z_10) );
  IV U4181 ( .A(n224), .Z(n2455) );
  AN2 U4182 ( .A(n2613), .B(n233), .Z(U3_U5_Z_1) );
  AN2 U4183 ( .A(n2613), .B(n234), .Z(U3_U5_Z_0) );
  AO4 U4184 ( .A(n2590), .B(n3851), .C(n3583), .D(n3852), .Z(U3_U4_Z_0) );
  ND2 U4185 ( .A(n3853), .B(n2197), .Z(n3852) );
  ND4 U4186 ( .A(n3854), .B(n3855), .C(n3856), .D(n3857), .Z(n3853) );
  NR4 U4187 ( .A(n4465), .B(n4469), .C(n4474), .D(n4479), .Z(n3857) );
  NR4 U4188 ( .A(n4484), .B(n4489), .C(n4494), .D(n4499), .Z(n3856) );
  NR4 U4189 ( .A(n4503), .B(n4507), .C(n4511), .D(n4515), .Z(n3855) );
  NR4 U4190 ( .A(n4519), .B(n4523), .C(n4527), .D(n4531), .Z(n3854) );
  ND2 U4191 ( .A(Datai[31]), .B(n3858), .Z(n3851) );
  ND4 U4192 ( .A(n3859), .B(n3860), .C(n3861), .D(n3862), .Z(n3858) );
  NR4 U4193 ( .A(Datai[9]), .B(Datai[8]), .C(Datai[7]), .D(Datai[6]), .Z(n3862) );
  NR4 U4194 ( .A(Datai[5]), .B(Datai[4]), .C(Datai[3]), .D(Datai[2]), .Z(n3861) );
  NR4 U4195 ( .A(Datai[1]), .B(Datai[15]), .C(Datai[14]), .D(Datai[13]), .Z(
        n3860) );
  NR4 U4196 ( .A(Datai[12]), .B(Datai[11]), .C(Datai[10]), .D(Datai[0]), .Z(
        n3859) );
  AO7 U4197 ( .A(n4569), .B(n3583), .C(n3863), .Z(U3_U3_Z_9) );
  AO7 U4198 ( .A(n4565), .B(n3583), .C(n3863), .Z(U3_U3_Z_8) );
  AO7 U4199 ( .A(n4561), .B(n3583), .C(n3863), .Z(U3_U3_Z_7) );
  EON1 U4200 ( .A(n2590), .B(n2745), .C(n4557), .D(n3864), .Z(U3_U3_Z_6) );
  IV U4201 ( .A(Datai[22]), .Z(n2745) );
  EON1 U4202 ( .A(n2590), .B(n2742), .C(n4553), .D(n3864), .Z(U3_U3_Z_5) );
  IV U4203 ( .A(Datai[21]), .Z(n2742) );
  EON1 U4204 ( .A(n2590), .B(n2739), .C(n4549), .D(n3864), .Z(U3_U3_Z_4) );
  IV U4205 ( .A(Datai[20]), .Z(n2739) );
  EON1 U4206 ( .A(n2590), .B(n2736), .C(n4545), .D(n3864), .Z(U3_U3_Z_3) );
  IV U4207 ( .A(Datai[19]), .Z(n2736) );
  EON1 U4208 ( .A(n2590), .B(n2733), .C(n4541), .D(n3864), .Z(U3_U3_Z_2) );
  IV U4209 ( .A(Datai[18]), .Z(n2733) );
  AO7 U4210 ( .A(n4589), .B(n3583), .C(n3863), .Z(U3_U3_Z_14) );
  AO7 U4211 ( .A(n4585), .B(n3583), .C(n3863), .Z(U3_U3_Z_13) );
  AO7 U4212 ( .A(n4581), .B(n3583), .C(n3863), .Z(U3_U3_Z_12) );
  AO7 U4213 ( .A(n4577), .B(n3583), .C(n3863), .Z(U3_U3_Z_11) );
  AO7 U4214 ( .A(n4573), .B(n3583), .C(n3863), .Z(U3_U3_Z_10) );
  ND2 U4215 ( .A(Datai[23]), .B(n2364), .Z(n3863) );
  IV U4216 ( .A(n2590), .Z(n2364) );
  EON1 U4217 ( .A(n2590), .B(n2730), .C(n4537), .D(n3864), .Z(U3_U3_Z_1) );
  IV U4218 ( .A(Datai[17]), .Z(n2730) );
  EON1 U4219 ( .A(n2590), .B(n2727), .C(n4533), .D(n3864), .Z(U3_U3_Z_0) );
  IV U4220 ( .A(Datai[16]), .Z(n2727) );
  NR2 U4221 ( .A(n3865), .B(n2154), .Z(U3_U2_Z_0) );
  AO2 U4222 ( .A(rEIP[0]), .B(n2246), .C(n2315), .D(rEIP[1]), .Z(n3865) );
  ND2 U4223 ( .A(n3866), .B(n2294), .Z(n2246) );
  IV U4224 ( .A(n3867), .Z(U3_U23_Z_0) );
  AO6 U4225 ( .A(n2550), .B(n3796), .C(n3815), .Z(n3867) );
  AO3 U4226 ( .A(n4505), .B(n3840), .C(n3868), .D(n3869), .Z(U3_U22_Z_9) );
  EO1 U4227 ( .A(n3870), .B(n4507), .C(n2357), .D(n4508), .Z(n3869) );
  ND2 U4228 ( .A(n3815), .B(n451), .Z(n3868) );
  AO3 U4229 ( .A(n4501), .B(n3840), .C(n3871), .D(n3872), .Z(U3_U22_Z_8) );
  EO1 U4230 ( .A(n3870), .B(n4503), .C(n2357), .D(n4504), .Z(n3872) );
  ND2 U4231 ( .A(n3815), .B(n452), .Z(n3871) );
  AO3 U4232 ( .A(n4496), .B(n3840), .C(n3873), .D(n3874), .Z(U3_U22_Z_7) );
  EO1 U4233 ( .A(n3870), .B(n4499), .C(n2357), .D(n4500), .Z(n3874) );
  ND2 U4234 ( .A(n3815), .B(n453), .Z(n3873) );
  AO3 U4235 ( .A(n4491), .B(n3840), .C(n3875), .D(n3876), .Z(U3_U22_Z_6) );
  EO1 U4236 ( .A(n3870), .B(n4494), .C(n2357), .D(n4495), .Z(n3876) );
  ND2 U4237 ( .A(n3815), .B(n454), .Z(n3875) );
  AO3 U4238 ( .A(n4486), .B(n3840), .C(n3877), .D(n3878), .Z(U3_U22_Z_5) );
  EO1 U4239 ( .A(n3870), .B(n4489), .C(n2357), .D(n4490), .Z(n3878) );
  ND2 U4240 ( .A(n3815), .B(n455), .Z(n3877) );
  AO3 U4241 ( .A(n4481), .B(n3840), .C(n3879), .D(n3880), .Z(U3_U22_Z_4) );
  EO1 U4242 ( .A(n3870), .B(n4484), .C(n2357), .D(n4485), .Z(n3880) );
  ND2 U4243 ( .A(n3815), .B(n456), .Z(n3879) );
  AO7 U4244 ( .A(n4646), .B(n3840), .C(n3824), .Z(U3_U22_Z_31) );
  AO4 U4245 ( .A(n3678), .B(n3824), .C(n4643), .D(n3840), .Z(U3_U22_Z_30) );
  IV U4246 ( .A(n430), .Z(n3678) );
  AO3 U4247 ( .A(n4476), .B(n3840), .C(n3881), .D(n3882), .Z(U3_U22_Z_3) );
  EO1 U4248 ( .A(n3870), .B(n4479), .C(n2357), .D(n4480), .Z(n3882) );
  ND2 U4249 ( .A(n3815), .B(n457), .Z(n3881) );
  AO4 U4250 ( .A(n3675), .B(n3824), .C(n4586), .D(n3840), .Z(U3_U22_Z_29) );
  IV U4251 ( .A(n431), .Z(n3675) );
  AO4 U4252 ( .A(n3672), .B(n3824), .C(n4582), .D(n3840), .Z(U3_U22_Z_28) );
  IV U4253 ( .A(n432), .Z(n3672) );
  AO4 U4254 ( .A(n3669), .B(n3824), .C(n4578), .D(n3840), .Z(U3_U22_Z_27) );
  IV U4255 ( .A(n433), .Z(n3669) );
  AO4 U4256 ( .A(n3666), .B(n3824), .C(n4574), .D(n3840), .Z(U3_U22_Z_26) );
  IV U4257 ( .A(n434), .Z(n3666) );
  AO4 U4258 ( .A(n3663), .B(n3824), .C(n4570), .D(n3840), .Z(U3_U22_Z_25) );
  IV U4259 ( .A(n435), .Z(n3663) );
  AO4 U4260 ( .A(n3660), .B(n3824), .C(n4566), .D(n3840), .Z(U3_U22_Z_24) );
  IV U4261 ( .A(n436), .Z(n3660) );
  AO7 U4262 ( .A(n3657), .B(n3824), .C(n3883), .Z(U3_U22_Z_23) );
  EO1 U4263 ( .A(n3826), .B(n3884), .C(n3840), .D(n4562), .Z(n3883) );
  AO7 U4264 ( .A(n2610), .B(n3885), .C(n3886), .Z(n3884) );
  EO1 U4265 ( .A(n3887), .B(n2145), .C(n3888), .D(n2570), .Z(n3886) );
  IV U4266 ( .A(n437), .Z(n3657) );
  AO3 U4267 ( .A(n3889), .B(n3812), .C(n3890), .D(n3891), .Z(U3_U22_Z_22) );
  AO2 U4268 ( .A(n3815), .B(n438), .C(n3892), .D(n3817), .Z(n3891) );
  OR2 U4269 ( .A(n3840), .B(n4558), .Z(n3890) );
  AO6 U4270 ( .A(n3893), .B(n3820), .C(n3894), .Z(n3889) );
  AO4 U4271 ( .A(n2570), .B(n3895), .C(n4468), .D(n3896), .Z(n3894) );
  AO3 U4272 ( .A(n3897), .B(n3812), .C(n3898), .D(n3899), .Z(U3_U22_Z_21) );
  AO2 U4273 ( .A(n3815), .B(n439), .C(n3900), .D(n3817), .Z(n3899) );
  OR2 U4274 ( .A(n3840), .B(n4554), .Z(n3898) );
  AO6 U4275 ( .A(n3901), .B(n3820), .C(n3902), .Z(n3897) );
  AO4 U4276 ( .A(n2570), .B(n3903), .C(n4468), .D(n3904), .Z(n3902) );
  AO3 U4277 ( .A(n3905), .B(n3812), .C(n3906), .D(n3907), .Z(U3_U22_Z_20) );
  AO2 U4278 ( .A(n3815), .B(n440), .C(n3908), .D(n3817), .Z(n3907) );
  OR2 U4279 ( .A(n3840), .B(n4550), .Z(n3906) );
  AO6 U4280 ( .A(n3909), .B(n3820), .C(n3910), .Z(n3905) );
  AO4 U4281 ( .A(n2570), .B(n3911), .C(n4468), .D(n3912), .Z(n3910) );
  AO3 U4282 ( .A(n4471), .B(n3840), .C(n3913), .D(n3914), .Z(U3_U22_Z_2) );
  EO1 U4283 ( .A(n3870), .B(n4474), .C(n2357), .D(n4475), .Z(n3914) );
  ND2 U4284 ( .A(n3815), .B(n458), .Z(n3913) );
  AO3 U4285 ( .A(n4529), .B(n3840), .C(n3915), .D(n3916), .Z(U3_U22_Z_15) );
  EO1 U4286 ( .A(n3870), .B(n4531), .C(n2357), .D(n4532), .Z(n3916) );
  ND2 U4287 ( .A(n3815), .B(n445), .Z(n3915) );
  AO3 U4288 ( .A(n4525), .B(n3840), .C(n3917), .D(n3918), .Z(U3_U22_Z_14) );
  EO1 U4289 ( .A(n3870), .B(n4527), .C(n2357), .D(n4528), .Z(n3918) );
  ND2 U4290 ( .A(n3815), .B(n446), .Z(n3917) );
  AO3 U4291 ( .A(n4521), .B(n3840), .C(n3919), .D(n3920), .Z(U3_U22_Z_13) );
  EO1 U4292 ( .A(n3870), .B(n4523), .C(n2357), .D(n4524), .Z(n3920) );
  ND2 U4293 ( .A(n3815), .B(n447), .Z(n3919) );
  AO3 U4294 ( .A(n4517), .B(n3840), .C(n3921), .D(n3922), .Z(U3_U22_Z_12) );
  EO1 U4295 ( .A(n3870), .B(n4519), .C(n2357), .D(n4520), .Z(n3922) );
  ND2 U4296 ( .A(n3815), .B(n448), .Z(n3921) );
  AO3 U4297 ( .A(n4513), .B(n3840), .C(n3923), .D(n3924), .Z(U3_U22_Z_11) );
  EO1 U4298 ( .A(n3870), .B(n4515), .C(n2357), .D(n4516), .Z(n3924) );
  ND2 U4299 ( .A(n3815), .B(n449), .Z(n3923) );
  AO3 U4300 ( .A(n4509), .B(n3840), .C(n3925), .D(n3926), .Z(U3_U22_Z_10) );
  EO1 U4301 ( .A(n3870), .B(n4511), .C(n2357), .D(n4512), .Z(n3926) );
  ND2 U4302 ( .A(n3815), .B(n450), .Z(n3925) );
  AO3 U4303 ( .A(n4452), .B(n3840), .C(n3927), .D(n3928), .Z(U3_U22_Z_1) );
  EO1 U4304 ( .A(n3870), .B(n4469), .C(n2357), .D(n4470), .Z(n3928) );
  ND2 U4305 ( .A(n3815), .B(n459), .Z(n3927) );
  AO3 U4306 ( .A(n4463), .B(n3840), .C(n3929), .D(n3930), .Z(U3_U22_Z_0) );
  EO1 U4307 ( .A(n3870), .B(n4465), .C(n2357), .D(n4466), .Z(n3930) );
  ND2 U4308 ( .A(n3815), .B(n460), .Z(n3929) );
  IV U4309 ( .A(n3824), .Z(n3815) );
  ND2 U4310 ( .A(n2389), .B(n2550), .Z(n3824) );
  AO6 U4311 ( .A(n2550), .B(n3796), .C(U3_U21_Z_0), .Z(n3840) );
  AO3 U4312 ( .A(n2598), .B(n2337), .C(n3931), .D(n3932), .Z(n2550) );
  OR3 U4313 ( .A(n4646), .B(n2245), .C(n2395), .Z(n3932) );
  ND2 U4314 ( .A(n4657), .B(n2581), .Z(n3931) );
  NR2 U4315 ( .A(n2261), .B(n4357), .Z(n2581) );
  IV U4316 ( .A(n2352), .Z(n2261) );
  AN3 U4317 ( .A(n2170), .B(n2151), .C(n2390), .Z(n2352) );
  IV U4318 ( .A(n429), .Z(n2337) );
  IV U4319 ( .A(n3933), .Z(U3_U21_Z_30) );
  AO1 U4320 ( .A(N1764), .B(n3870), .C(n3934), .D(n3935), .Z(n3933) );
  AO7 U4321 ( .A(n3936), .B(n2228), .C(n3937), .Z(n3935) );
  AO2 U4322 ( .A(n4633), .B(n3938), .C(n3887), .D(n3939), .Z(n3937) );
  AO4 U4323 ( .A(n2167), .B(n3940), .C(n3941), .D(n3942), .Z(n3887) );
  AO4 U4324 ( .A(n4634), .B(n3943), .C(n3944), .D(n3945), .Z(n3942) );
  AN2 U4325 ( .A(n2167), .B(n4378), .Z(n3944) );
  NR2 U4326 ( .A(n4376), .B(n2349), .Z(n3941) );
  AO4 U4327 ( .A(n3888), .B(n3946), .C(n2357), .D(n4642), .Z(n3934) );
  IV U4328 ( .A(n3947), .Z(U3_U21_Z_29) );
  AO1 U4329 ( .A(N1763), .B(n3870), .C(n3948), .D(n3949), .Z(n3947) );
  ND2 U4330 ( .A(n3950), .B(n3951), .Z(n3949) );
  EO1 U4331 ( .A(n4391), .B(n3952), .C(n3896), .D(n3953), .Z(n3951) );
  AO3 U4332 ( .A(n4629), .B(n3943), .C(n2167), .D(n3954), .Z(n3896) );
  IV U4333 ( .A(n3955), .Z(n3954) );
  AO4 U4334 ( .A(n2349), .B(n4387), .C(n2347), .D(n4625), .Z(n3955) );
  AO2 U4335 ( .A(n3892), .B(n3956), .C(n4628), .D(n3957), .Z(n3950) );
  AO4 U4336 ( .A(n3895), .B(n3946), .C(n2357), .D(n4641), .Z(n3948) );
  IV U4337 ( .A(n3958), .Z(U3_U21_Z_28) );
  AO1 U4338 ( .A(N1762), .B(n3870), .C(n3959), .D(n3960), .Z(n3958) );
  AO3 U4339 ( .A(n3953), .B(n3904), .C(n3961), .D(n3962), .Z(n3960) );
  ND2 U4340 ( .A(n3900), .B(n3956), .Z(n3962) );
  AO2 U4341 ( .A(n4370), .B(n3952), .C(n4621), .D(n3938), .Z(n3961) );
  AO3 U4342 ( .A(n4622), .B(n3943), .C(n2167), .D(n3963), .Z(n3904) );
  IV U4343 ( .A(n3964), .Z(n3963) );
  AO4 U4344 ( .A(n2349), .B(n4366), .C(n2347), .D(n4619), .Z(n3964) );
  AO4 U4345 ( .A(n3903), .B(n3946), .C(n2357), .D(n4640), .Z(n3959) );
  IV U4346 ( .A(n3965), .Z(U3_U21_Z_27) );
  AO1 U4347 ( .A(N1761), .B(n3870), .C(n3966), .D(n3967), .Z(n3965) );
  AO3 U4348 ( .A(n3953), .B(n3912), .C(n3968), .D(n3969), .Z(n3967) );
  ND2 U4349 ( .A(n3908), .B(n3956), .Z(n3969) );
  AO2 U4350 ( .A(n4444), .B(n3952), .C(n4615), .D(n3938), .Z(n3968) );
  AO3 U4351 ( .A(n4616), .B(n3943), .C(n2167), .D(n3970), .Z(n3912) );
  IV U4352 ( .A(n3971), .Z(n3970) );
  AO4 U4353 ( .A(n2349), .B(n4440), .C(n2347), .D(n4613), .Z(n3971) );
  AO4 U4354 ( .A(n3911), .B(n3946), .C(n2357), .D(n4639), .Z(n3966) );
  IV U4355 ( .A(n3972), .Z(U3_U21_Z_26) );
  AO1 U4356 ( .A(N1760), .B(n3870), .C(n3973), .D(n3974), .Z(n3972) );
  AO3 U4357 ( .A(n3953), .B(n3823), .C(n3975), .D(n3976), .Z(n3974) );
  ND2 U4358 ( .A(n3816), .B(n3956), .Z(n3976) );
  NR2 U4359 ( .A(n3953), .B(n2167), .Z(n3956) );
  AO2 U4360 ( .A(n4434), .B(n3952), .C(n4609), .D(n3938), .Z(n3975) );
  AO3 U4361 ( .A(n4610), .B(n3943), .C(n2167), .D(n3977), .Z(n3823) );
  IV U4362 ( .A(n3978), .Z(n3977) );
  AO4 U4363 ( .A(n2349), .B(n4430), .C(n2347), .D(n4607), .Z(n3978) );
  IV U4364 ( .A(n3939), .Z(n3953) );
  AO4 U4365 ( .A(n3946), .B(n3822), .C(n2357), .D(n4638), .Z(n3973) );
  IV U4366 ( .A(n3979), .Z(U3_U21_Z_25) );
  AO1 U4367 ( .A(N1759), .B(n3870), .C(n3980), .D(n3981), .Z(n3979) );
  AO7 U4368 ( .A(n3936), .B(n2229), .C(n3982), .Z(n3981) );
  AO2 U4369 ( .A(n3830), .B(n3939), .C(n4603), .D(n3957), .Z(n3982) );
  AO4 U4370 ( .A(n2167), .B(n3983), .C(n3984), .D(n3985), .Z(n3830) );
  AO4 U4371 ( .A(n4604), .B(n3943), .C(n3986), .D(n3945), .Z(n3985) );
  AN2 U4372 ( .A(n2167), .B(n4398), .Z(n3986) );
  NR2 U4373 ( .A(n4396), .B(n2349), .Z(n3984) );
  AO4 U4374 ( .A(n3831), .B(n3946), .C(n2357), .D(n4637), .Z(n3980) );
  IV U4375 ( .A(n3987), .Z(U3_U21_Z_24) );
  AO1 U4376 ( .A(N1758), .B(n3870), .C(n3988), .D(n3989), .Z(n3987) );
  AO7 U4377 ( .A(n3936), .B(n2230), .C(n3990), .Z(n3989) );
  AO2 U4378 ( .A(n4597), .B(n3938), .C(n3836), .D(n3939), .Z(n3990) );
  AO4 U4379 ( .A(n2167), .B(n3991), .C(n3992), .D(n3993), .Z(n3836) );
  AO4 U4380 ( .A(n4598), .B(n3943), .C(n3994), .D(n3945), .Z(n3993) );
  AN2 U4381 ( .A(n2167), .B(n4420), .Z(n3994) );
  NR2 U4382 ( .A(n4418), .B(n2349), .Z(n3992) );
  AO4 U4383 ( .A(n3837), .B(n3946), .C(n2357), .D(n4636), .Z(n3988) );
  IV U4384 ( .A(n3817), .Z(n3946) );
  AO3 U4385 ( .A(n2265), .B(n3795), .C(n3995), .D(n3996), .Z(U3_U21_Z_23) );
  AO6 U4386 ( .A(n3939), .B(n3843), .C(n3997), .Z(n3996) );
  IV U4387 ( .A(n3998), .Z(n3997) );
  AO2 U4388 ( .A(n4411), .B(n3952), .C(n4592), .D(n3938), .Z(n3998) );
  NR2 U4389 ( .A(n3999), .B(n3943), .Z(n3938) );
  IV U4390 ( .A(n3936), .Z(n3952) );
  ND2 U4391 ( .A(n3957), .B(n4000), .Z(n3936) );
  IV U4392 ( .A(n3999), .Z(n3957) );
  ND2 U4393 ( .A(n3826), .B(n2578), .Z(n3999) );
  AO4 U4394 ( .A(n2167), .B(n4001), .C(n4002), .D(n4003), .Z(n3843) );
  AO4 U4395 ( .A(n4593), .B(n3943), .C(n4004), .D(n3945), .Z(n4003) );
  NR2 U4396 ( .A(n4000), .B(n4461), .Z(n3945) );
  AN2 U4397 ( .A(n2167), .B(n4408), .Z(n4004) );
  NR2 U4398 ( .A(n4406), .B(n2349), .Z(n4002) );
  NR2 U4399 ( .A(n3812), .B(n2145), .Z(n3939) );
  EO1 U4400 ( .A(n3844), .B(n3817), .C(n2357), .D(n4631), .Z(n3995) );
  NR2 U4401 ( .A(n3812), .B(n4005), .Z(n3817) );
  IV U4402 ( .A(N1757), .Z(n2265) );
  AO4 U4403 ( .A(n2894), .B(n3795), .C(n4624), .D(n2357), .Z(U3_U21_Z_22) );
  IV U4404 ( .A(N1756), .Z(n2894) );
  AO4 U4405 ( .A(n2890), .B(n3795), .C(n4618), .D(n2357), .Z(U3_U21_Z_21) );
  IV U4406 ( .A(N1755), .Z(n2890) );
  AO4 U4407 ( .A(n2886), .B(n3795), .C(n4612), .D(n2357), .Z(U3_U21_Z_20) );
  IV U4408 ( .A(N1754), .Z(n2886) );
  AO4 U4409 ( .A(n2882), .B(n3795), .C(n4606), .D(n2357), .Z(U3_U21_Z_19) );
  IV U4410 ( .A(N1753), .Z(n2882) );
  AO4 U4411 ( .A(n2878), .B(n3795), .C(n4600), .D(n2357), .Z(U3_U21_Z_18) );
  IV U4412 ( .A(N1752), .Z(n2878) );
  AO4 U4413 ( .A(n2874), .B(n3795), .C(n4595), .D(n2357), .Z(U3_U21_Z_17) );
  IV U4414 ( .A(N1751), .Z(n2874) );
  AO4 U4415 ( .A(n2867), .B(n3795), .C(n4590), .D(n2357), .Z(U3_U21_Z_16) );
  ND3 U4416 ( .A(n2170), .B(n4658), .C(n2390), .Z(n2357) );
  IV U4417 ( .A(N1750), .Z(n2867) );
  NR2 U4418 ( .A(n2726), .B(n2359), .Z(U3_U21_Z_0) );
  ND2 U4419 ( .A(n4006), .B(n4007), .Z(n2726) );
  AO4 U4420 ( .A(n2166), .B(n3866), .C(n2191), .D(n2294), .Z(U3_U1_Z_9) );
  AO4 U4421 ( .A(n2191), .B(n3866), .C(n2163), .D(n2294), .Z(U3_U1_Z_8) );
  AO4 U4422 ( .A(n2163), .B(n3866), .C(n2192), .D(n2294), .Z(U3_U1_Z_7) );
  AO4 U4423 ( .A(n2192), .B(n3866), .C(n2152), .D(n2294), .Z(U3_U1_Z_6) );
  AO4 U4424 ( .A(n2152), .B(n3866), .C(n2172), .D(n2294), .Z(U3_U1_Z_5) );
  AO4 U4425 ( .A(n2172), .B(n3866), .C(n2153), .D(n2294), .Z(U3_U1_Z_4) );
  AO4 U4426 ( .A(n2153), .B(n3866), .C(n2173), .D(n2294), .Z(U3_U1_Z_3) );
  AO4 U4427 ( .A(n2154), .B(n3866), .C(n2174), .D(n2294), .Z(U3_U1_Z_29) );
  AO4 U4428 ( .A(n2174), .B(n3866), .C(n2156), .D(n2294), .Z(U3_U1_Z_28) );
  AO4 U4429 ( .A(n2156), .B(n3866), .C(n2175), .D(n2294), .Z(U3_U1_Z_27) );
  AO4 U4430 ( .A(n2175), .B(n3866), .C(n2157), .D(n2294), .Z(U3_U1_Z_26) );
  AO4 U4431 ( .A(n2157), .B(n3866), .C(n2176), .D(n2294), .Z(U3_U1_Z_25) );
  AO4 U4432 ( .A(n2176), .B(n3866), .C(n2158), .D(n2294), .Z(U3_U1_Z_24) );
  AO4 U4433 ( .A(n2158), .B(n3866), .C(n2177), .D(n2294), .Z(U3_U1_Z_23) );
  AO4 U4434 ( .A(n2177), .B(n3866), .C(n2159), .D(n2294), .Z(U3_U1_Z_22) );
  AO4 U4435 ( .A(n2159), .B(n3866), .C(n2178), .D(n2294), .Z(U3_U1_Z_21) );
  AO4 U4436 ( .A(n2178), .B(n3866), .C(n2160), .D(n2294), .Z(U3_U1_Z_20) );
  AO4 U4437 ( .A(n2173), .B(n3866), .C(n2155), .D(n2294), .Z(U3_U1_Z_2) );
  AO4 U4438 ( .A(n2160), .B(n3866), .C(n2179), .D(n2294), .Z(U3_U1_Z_19) );
  AO4 U4439 ( .A(n2179), .B(n3866), .C(n2161), .D(n2294), .Z(U3_U1_Z_18) );
  AO4 U4440 ( .A(n2161), .B(n3866), .C(n2181), .D(n2294), .Z(U3_U1_Z_17) );
  AO4 U4441 ( .A(n2181), .B(n3866), .C(n2162), .D(n2294), .Z(U3_U1_Z_16) );
  AO4 U4442 ( .A(n2162), .B(n3866), .C(n2182), .D(n2294), .Z(U3_U1_Z_15) );
  AO4 U4443 ( .A(n2182), .B(n3866), .C(n2164), .D(n2294), .Z(U3_U1_Z_14) );
  AO4 U4444 ( .A(n2164), .B(n3866), .C(n2193), .D(n2294), .Z(U3_U1_Z_13) );
  AO4 U4445 ( .A(n2193), .B(n3866), .C(n2165), .D(n2294), .Z(U3_U1_Z_12) );
  AO4 U4446 ( .A(n2165), .B(n3866), .C(n2194), .D(n2294), .Z(U3_U1_Z_11) );
  AO4 U4447 ( .A(n2194), .B(n3866), .C(n2166), .D(n2294), .Z(U3_U1_Z_10) );
  AO4 U4448 ( .A(n2155), .B(n3866), .C(n2180), .D(n2294), .Z(U3_U1_Z_1) );
  AO4 U4449 ( .A(n2180), .B(n3866), .C(n2149), .D(n2294), .Z(U3_U1_Z_0) );
  ND2 U4450 ( .A(n2308), .B(n2212), .Z(n2294) );
  NR2 U4451 ( .A(n4651), .B(n4667), .Z(n2308) );
  IV U4452 ( .A(n2315), .Z(n3866) );
  AO3 U4453 ( .A(n4008), .B(n2231), .C(n4009), .D(n4010), .Z(U3_U19_Z_7) );
  ND2 U4454 ( .A(n4011), .B(n2253), .Z(n4009) );
  AO3 U4455 ( .A(n4008), .B(n2232), .C(n4012), .D(n4010), .Z(U3_U19_Z_6) );
  ND2 U4456 ( .A(n4013), .B(n2253), .Z(n4012) );
  IV U4457 ( .A(n4014), .Z(n4013) );
  AO3 U4458 ( .A(n4008), .B(n2233), .C(n4015), .D(n4010), .Z(U3_U19_Z_5) );
  ND2 U4459 ( .A(n4016), .B(n2253), .Z(n4015) );
  IV U4460 ( .A(n4017), .Z(n4016) );
  AO3 U4461 ( .A(n4008), .B(n2234), .C(n4018), .D(n4010), .Z(U3_U19_Z_4) );
  ND2 U4462 ( .A(n4019), .B(n2253), .Z(n4018) );
  IV U4463 ( .A(n4020), .Z(n4019) );
  AO3 U4464 ( .A(n4008), .B(n2235), .C(n4021), .D(n4010), .Z(U3_U19_Z_3) );
  ND2 U4465 ( .A(n4022), .B(n2253), .Z(n4021) );
  IV U4466 ( .A(n4023), .Z(n4022) );
  AO3 U4467 ( .A(n4008), .B(n2236), .C(n4024), .D(n4010), .Z(U3_U19_Z_2) );
  ND2 U4468 ( .A(n4025), .B(n2253), .Z(n4024) );
  IV U4469 ( .A(n4026), .Z(n4025) );
  AO3 U4470 ( .A(n2372), .B(n4027), .C(n4010), .D(n4028), .Z(U3_U19_Z_0) );
  AO2 U4471 ( .A(n4029), .B(n2253), .C(n4413), .D(n2254), .Z(n4028) );
  OR3 U4472 ( .A(n4030), .B(n3810), .C(n4031), .Z(n2253) );
  IV U4473 ( .A(n4032), .Z(n4029) );
  ND2 U4474 ( .A(n2250), .B(n2387), .Z(n4027) );
  ND3 U4475 ( .A(n4033), .B(n4034), .C(n4035), .Z(n2250) );
  AO3 U4476 ( .A(n4358), .B(n3690), .C(n4036), .D(n4037), .Z(U3_U18_Z_9) );
  AO2 U4477 ( .A(n451), .B(n4038), .C(rEIP[9]), .D(n2251), .Z(n4037) );
  AO7 U4478 ( .A(n4039), .B(n4040), .C(n2613), .Z(n4036) );
  AO4 U4479 ( .A(n4005), .B(n3834), .C(n2610), .D(n4041), .Z(n4040) );
  AO4 U4480 ( .A(n2570), .B(n3991), .C(n2348), .D(n3837), .Z(n4039) );
  AO7 U4481 ( .A(n4429), .B(n2347), .C(n4042), .Z(n3837) );
  IV U4482 ( .A(n4043), .Z(n4042) );
  AO4 U4483 ( .A(n3943), .B(n4599), .C(n2349), .D(n4427), .Z(n4043) );
  AO3 U4484 ( .A(n4359), .B(n3690), .C(n4044), .D(n4045), .Z(U3_U18_Z_8) );
  AO2 U4485 ( .A(n452), .B(n4038), .C(rEIP[8]), .D(n2251), .Z(n4045) );
  AO7 U4486 ( .A(n4046), .B(n4047), .C(n2613), .Z(n4044) );
  AO4 U4487 ( .A(n4005), .B(n3841), .C(n2610), .D(n4048), .Z(n4047) );
  EON1 U4488 ( .A(n2570), .B(n4001), .C(n2578), .D(n3844), .Z(n4046) );
  AO6 U4489 ( .A(n2237), .B(n4000), .C(n4049), .Z(n3844) );
  AO4 U4490 ( .A(n3943), .B(n4594), .C(n2349), .D(n4415), .Z(n4049) );
  AO7 U4491 ( .A(n2368), .B(n2152), .C(n4050), .Z(U3_U18_Z_7) );
  AO2 U4492 ( .A(n4498), .B(n4051), .C(n453), .D(n4038), .Z(n4050) );
  AO7 U4493 ( .A(n2368), .B(n2172), .C(n4052), .Z(U3_U18_Z_6) );
  AO2 U4494 ( .A(n4493), .B(n4051), .C(n454), .D(n4038), .Z(n4052) );
  AO7 U4495 ( .A(n2368), .B(n2153), .C(n4053), .Z(U3_U18_Z_5) );
  AO2 U4496 ( .A(n4488), .B(n4051), .C(n455), .D(n4038), .Z(n4053) );
  AO7 U4497 ( .A(n2368), .B(n2173), .C(n4054), .Z(U3_U18_Z_4) );
  AO2 U4498 ( .A(n4483), .B(n4051), .C(n456), .D(n4038), .Z(n4054) );
  AO7 U4499 ( .A(n2368), .B(n2154), .C(n4055), .Z(U3_U18_Z_31) );
  AO2 U4500 ( .A(n4657), .B(n4051), .C(n429), .D(n4038), .Z(n4055) );
  AO7 U4501 ( .A(n2368), .B(n2174), .C(n4056), .Z(U3_U18_Z_30) );
  AO2 U4502 ( .A(n4645), .B(n4051), .C(n430), .D(n4038), .Z(n4056) );
  AO7 U4503 ( .A(n2368), .B(n2155), .C(n4057), .Z(U3_U18_Z_3) );
  AO2 U4504 ( .A(n4478), .B(n4051), .C(n457), .D(n4038), .Z(n4057) );
  AO7 U4505 ( .A(n2368), .B(n2156), .C(n4058), .Z(U3_U18_Z_29) );
  AO2 U4506 ( .A(n4588), .B(n4051), .C(n431), .D(n4038), .Z(n4058) );
  AO7 U4507 ( .A(n2368), .B(n2175), .C(n4059), .Z(U3_U18_Z_28) );
  AO2 U4508 ( .A(n4584), .B(n4051), .C(n432), .D(n4038), .Z(n4059) );
  AO7 U4509 ( .A(n2368), .B(n2157), .C(n4060), .Z(U3_U18_Z_27) );
  AO2 U4510 ( .A(n4580), .B(n4051), .C(n433), .D(n4038), .Z(n4060) );
  AO7 U4511 ( .A(n2368), .B(n2176), .C(n4061), .Z(U3_U18_Z_26) );
  AO2 U4512 ( .A(n4576), .B(n4051), .C(n434), .D(n4038), .Z(n4061) );
  AO7 U4513 ( .A(n2368), .B(n2158), .C(n4062), .Z(U3_U18_Z_25) );
  AO2 U4514 ( .A(n4572), .B(n4051), .C(n435), .D(n4038), .Z(n4062) );
  AO7 U4515 ( .A(n2368), .B(n2177), .C(n4063), .Z(U3_U18_Z_24) );
  AO2 U4516 ( .A(n4568), .B(n4051), .C(n436), .D(n4038), .Z(n4063) );
  AO7 U4517 ( .A(n2368), .B(n2159), .C(n4064), .Z(U3_U18_Z_23) );
  AO2 U4518 ( .A(n4564), .B(n4051), .C(n437), .D(n4038), .Z(n4064) );
  AO7 U4519 ( .A(n2368), .B(n2178), .C(n4065), .Z(U3_U18_Z_22) );
  AO2 U4520 ( .A(n4560), .B(n4051), .C(n438), .D(n4038), .Z(n4065) );
  AO7 U4521 ( .A(n2368), .B(n2160), .C(n4066), .Z(U3_U18_Z_21) );
  AO2 U4522 ( .A(n4556), .B(n4051), .C(n439), .D(n4038), .Z(n4066) );
  AO7 U4523 ( .A(n2368), .B(n2179), .C(n4067), .Z(U3_U18_Z_20) );
  AO2 U4524 ( .A(n4552), .B(n4051), .C(n440), .D(n4038), .Z(n4067) );
  AO7 U4525 ( .A(n2368), .B(n2180), .C(n4068), .Z(U3_U18_Z_2) );
  AO2 U4526 ( .A(n4473), .B(n4051), .C(n458), .D(n4038), .Z(n4068) );
  AO7 U4527 ( .A(n2368), .B(n2161), .C(n4069), .Z(U3_U18_Z_19) );
  AO2 U4528 ( .A(n4548), .B(n4051), .C(n441), .D(n4038), .Z(n4069) );
  AO7 U4529 ( .A(n2368), .B(n2181), .C(n4070), .Z(U3_U18_Z_18) );
  AO2 U4530 ( .A(n4544), .B(n4051), .C(n442), .D(n4038), .Z(n4070) );
  AO7 U4531 ( .A(n2368), .B(n2162), .C(n4071), .Z(U3_U18_Z_17) );
  AO2 U4532 ( .A(n4540), .B(n4051), .C(n443), .D(n4038), .Z(n4071) );
  AO7 U4533 ( .A(n2368), .B(n2182), .C(n4072), .Z(U3_U18_Z_16) );
  AO2 U4534 ( .A(n4536), .B(n4051), .C(n444), .D(n4038), .Z(n4072) );
  AO3 U4535 ( .A(n4360), .B(n3690), .C(n4073), .D(n4074), .Z(U3_U18_Z_15) );
  AO2 U4536 ( .A(n445), .B(n4038), .C(rEIP[15]), .D(n2251), .Z(n4074) );
  AO7 U4537 ( .A(n4075), .B(n4076), .C(n2613), .Z(n4073) );
  EON1 U4538 ( .A(n4005), .B(n3885), .C(n3820), .D(n4077), .Z(n4076) );
  AO4 U4539 ( .A(n2570), .B(n3940), .C(n2348), .D(n3888), .Z(n4075) );
  AO7 U4540 ( .A(n4386), .B(n2347), .C(n4078), .Z(n3888) );
  IV U4541 ( .A(n4079), .Z(n4078) );
  AO4 U4542 ( .A(n3943), .B(n4635), .C(n2349), .D(n4384), .Z(n4079) );
  AO3 U4543 ( .A(n4361), .B(n3690), .C(n4080), .D(n4081), .Z(U3_U18_Z_14) );
  AO2 U4544 ( .A(n446), .B(n4038), .C(rEIP[14]), .D(n2251), .Z(n4081) );
  AO7 U4545 ( .A(n4082), .B(n4083), .C(n2613), .Z(n4080) );
  AO4 U4546 ( .A(n4005), .B(n4084), .C(n2610), .D(n4085), .Z(n4083) );
  EON1 U4547 ( .A(n2348), .B(n3895), .C(n2573), .D(n3892), .Z(n4082) );
  AO7 U4548 ( .A(n4626), .B(n2347), .C(n4086), .Z(n3895) );
  IV U4549 ( .A(n4087), .Z(n4086) );
  AO4 U4550 ( .A(n3943), .B(n4630), .C(n2349), .D(n4394), .Z(n4087) );
  AO3 U4551 ( .A(n4362), .B(n3690), .C(n4088), .D(n4089), .Z(U3_U18_Z_13) );
  AO2 U4552 ( .A(n447), .B(n4038), .C(rEIP[13]), .D(n2251), .Z(n4089) );
  AO7 U4553 ( .A(n4090), .B(n4091), .C(n2613), .Z(n4088) );
  AO4 U4554 ( .A(n4005), .B(n4092), .C(n2610), .D(n4093), .Z(n4091) );
  EON1 U4555 ( .A(n2348), .B(n3903), .C(n2573), .D(n3900), .Z(n4090) );
  AO7 U4556 ( .A(n4375), .B(n2347), .C(n4094), .Z(n3903) );
  IV U4557 ( .A(n4095), .Z(n4094) );
  AO4 U4558 ( .A(n3943), .B(n4623), .C(n2349), .D(n4373), .Z(n4095) );
  AO3 U4559 ( .A(n4363), .B(n3690), .C(n4096), .D(n4097), .Z(U3_U18_Z_12) );
  AO2 U4560 ( .A(n448), .B(n4038), .C(rEIP[12]), .D(n2251), .Z(n4097) );
  AO7 U4561 ( .A(n4098), .B(n4099), .C(n2613), .Z(n4096) );
  AO4 U4562 ( .A(n4005), .B(n4100), .C(n2610), .D(n4101), .Z(n4099) );
  EON1 U4563 ( .A(n2348), .B(n3911), .C(n2573), .D(n3908), .Z(n4098) );
  AO7 U4564 ( .A(n4449), .B(n2347), .C(n4102), .Z(n3911) );
  IV U4565 ( .A(n4103), .Z(n4102) );
  AO4 U4566 ( .A(n3943), .B(n4617), .C(n2349), .D(n4447), .Z(n4103) );
  AO3 U4567 ( .A(n4364), .B(n3690), .C(n4104), .D(n4105), .Z(U3_U18_Z_11) );
  AO2 U4568 ( .A(n449), .B(n4038), .C(rEIP[11]), .D(n2251), .Z(n4105) );
  AO7 U4569 ( .A(n4106), .B(n4107), .C(n2613), .Z(n4104) );
  AO4 U4570 ( .A(n4005), .B(n4108), .C(n2610), .D(n4109), .Z(n4107) );
  EON1 U4571 ( .A(n2348), .B(n3822), .C(n2573), .D(n3816), .Z(n4106) );
  AO7 U4572 ( .A(n4439), .B(n2347), .C(n4110), .Z(n3822) );
  IV U4573 ( .A(n4111), .Z(n4110) );
  AO4 U4574 ( .A(n3943), .B(n4611), .C(n2349), .D(n4437), .Z(n4111) );
  AO3 U4575 ( .A(n4365), .B(n3690), .C(n4112), .D(n4113), .Z(U3_U18_Z_10) );
  AO2 U4576 ( .A(n450), .B(n4038), .C(rEIP[10]), .D(n2251), .Z(n4113) );
  AO7 U4577 ( .A(n4114), .B(n4115), .C(n2613), .Z(n4112) );
  AO4 U4578 ( .A(n4005), .B(n3828), .C(n2610), .D(n4116), .Z(n4115) );
  AO4 U4579 ( .A(n2570), .B(n3983), .C(n2348), .D(n3831), .Z(n4114) );
  AO7 U4580 ( .A(n4601), .B(n2347), .C(n4117), .Z(n3831) );
  IV U4581 ( .A(n4118), .Z(n4117) );
  AO4 U4582 ( .A(n3943), .B(n4605), .C(n2349), .D(n4404), .Z(n4118) );
  IV U4583 ( .A(n4051), .Z(n3690) );
  AO7 U4584 ( .A(n2368), .B(n2149), .C(n4119), .Z(U3_U18_Z_1) );
  AO2 U4585 ( .A(n4453), .B(n4051), .C(n459), .D(n4038), .Z(n4119) );
  AO7 U4586 ( .A(n2368), .B(n2168), .C(n4120), .Z(U3_U18_Z_0) );
  AO2 U4587 ( .A(n4654), .B(n4051), .C(n460), .D(n4038), .Z(n4120) );
  OR3 U4588 ( .A(n3810), .B(U3_U14_Z_7), .C(n4030), .Z(n4038) );
  AO7 U4589 ( .A(n3586), .B(n2372), .C(n2248), .Z(n4051) );
  AO6 U4590 ( .A(n3691), .B(n4121), .C(n2779), .Z(n2248) );
  ND2 U4591 ( .A(n3582), .B(n4122), .Z(n2779) );
  ND3 U4592 ( .A(n3805), .B(n2286), .C(n2392), .Z(n4122) );
  IV U4593 ( .A(n3808), .Z(n2392) );
  IV U4594 ( .A(n2283), .Z(n4121) );
  AN3 U4595 ( .A(n2284), .B(n2286), .C(n3805), .Z(n3691) );
  IV U4596 ( .A(n2251), .Z(n2368) );
  AN3 U4597 ( .A(n2288), .B(n3805), .C(n2548), .Z(n2251) );
  NR2 U4598 ( .A(n2553), .B(n2287), .Z(n2548) );
  ND2 U4599 ( .A(n4665), .B(n2286), .Z(n2553) );
  NR2 U4600 ( .A(n4014), .B(n4010), .Z(U3_U14_Z_6) );
  AO3 U4601 ( .A(n3892), .B(n2348), .C(n4123), .D(n4124), .Z(n4014) );
  AO2 U4602 ( .A(n2573), .B(n4084), .C(n3820), .D(n4125), .Z(n4124) );
  ND2 U4603 ( .A(n2571), .B(n4085), .Z(n4123) );
  IV U4604 ( .A(n4126), .Z(n4085) );
  AO6 U4605 ( .A(n2238), .B(n4000), .C(n4127), .Z(n3892) );
  AO4 U4606 ( .A(n3943), .B(n4392), .C(n2349), .D(n4393), .Z(n4127) );
  NR2 U4607 ( .A(n4017), .B(n4010), .Z(U3_U14_Z_5) );
  AO3 U4608 ( .A(n3900), .B(n2348), .C(n4128), .D(n4129), .Z(n4017) );
  MUX21L U4609 ( .A(n4092), .B(n4130), .S(n4461), .Z(n4129) );
  ND2 U4610 ( .A(n2571), .B(n4093), .Z(n4128) );
  IV U4611 ( .A(n4131), .Z(n4093) );
  AO6 U4612 ( .A(n2239), .B(n4000), .C(n4132), .Z(n3900) );
  AO4 U4613 ( .A(n3943), .B(n4371), .C(n2349), .D(n4372), .Z(n4132) );
  NR2 U4614 ( .A(n4020), .B(n4010), .Z(U3_U14_Z_4) );
  AO3 U4615 ( .A(n3908), .B(n2348), .C(n4133), .D(n4134), .Z(n4020) );
  AO2 U4616 ( .A(n2573), .B(n4100), .C(n3820), .D(n4135), .Z(n4134) );
  ND2 U4617 ( .A(n2571), .B(n4101), .Z(n4133) );
  IV U4618 ( .A(n4136), .Z(n4101) );
  AO6 U4619 ( .A(n2240), .B(n4000), .C(n4137), .Z(n3908) );
  AO4 U4620 ( .A(n3943), .B(n4445), .C(n2349), .D(n4446), .Z(n4137) );
  NR2 U4621 ( .A(n4023), .B(n4010), .Z(U3_U14_Z_3) );
  AO3 U4622 ( .A(n3816), .B(n2348), .C(n4138), .D(n4139), .Z(n4023) );
  MUX21L U4623 ( .A(n4108), .B(n4140), .S(n4461), .Z(n4139) );
  ND2 U4624 ( .A(n2571), .B(n4109), .Z(n4138) );
  IV U4625 ( .A(n4141), .Z(n4109) );
  AO6 U4626 ( .A(n2241), .B(n4000), .C(n4142), .Z(n3816) );
  AO4 U4627 ( .A(n3943), .B(n4435), .C(n2349), .D(n4436), .Z(n4142) );
  IV U4628 ( .A(n2347), .Z(n4000) );
  AO3 U4629 ( .A(n4026), .B(n4010), .C(n2590), .D(n4143), .Z(U3_U14_Z_2) );
  ND2 U4630 ( .A(n4144), .B(n4145), .Z(n4026) );
  AO2 U4631 ( .A(n2578), .B(n3983), .C(n2571), .D(n4116), .Z(n4145) );
  IV U4632 ( .A(n4146), .Z(n4116) );
  AO7 U4633 ( .A(n4602), .B(n2347), .C(n4147), .Z(n3983) );
  IV U4634 ( .A(n4148), .Z(n4147) );
  AO4 U4635 ( .A(n3943), .B(n4402), .C(n2349), .D(n4403), .Z(n4148) );
  AO2 U4636 ( .A(n2573), .B(n3828), .C(n3820), .D(n4149), .Z(n4144) );
  IV U4637 ( .A(n4150), .Z(U3_U14_Z_1) );
  AO1 U4638 ( .A(n2252), .B(U3_U14_Z_7), .C(n4151), .D(n4152), .Z(n4150) );
  ND2 U4639 ( .A(n4153), .B(n3540), .Z(n4152) );
  AN2 U4640 ( .A(n4154), .B(n4155), .Z(n2252) );
  AO2 U4641 ( .A(n2578), .B(n3991), .C(n2571), .D(n4041), .Z(n4155) );
  IV U4642 ( .A(n4156), .Z(n4041) );
  AO7 U4643 ( .A(n4596), .B(n2347), .C(n4157), .Z(n3991) );
  IV U4644 ( .A(n4158), .Z(n4157) );
  AO4 U4645 ( .A(n3943), .B(n4424), .C(n2349), .D(n4426), .Z(n4158) );
  AO2 U4646 ( .A(n2573), .B(n3834), .C(n3820), .D(n4159), .Z(n4154) );
  AO3 U4647 ( .A(n4032), .B(n4010), .C(n2778), .D(n4143), .Z(U3_U14_Z_0) );
  IV U4648 ( .A(n4160), .Z(n2778) );
  ND2 U4649 ( .A(n4161), .B(n4162), .Z(n4032) );
  AO2 U4650 ( .A(n2578), .B(n4001), .C(n2571), .D(n4048), .Z(n4162) );
  IV U4651 ( .A(n4163), .Z(n4048) );
  AO7 U4652 ( .A(n4591), .B(n2347), .C(n4164), .Z(n4001) );
  IV U4653 ( .A(n4165), .Z(n4164) );
  AO4 U4654 ( .A(n3943), .B(n4412), .C(n2349), .D(n4414), .Z(n4165) );
  AO2 U4655 ( .A(n2573), .B(n3841), .C(n3820), .D(n4166), .Z(n4161) );
  IV U4656 ( .A(n2570), .Z(n2573) );
  AO3 U4657 ( .A(n4506), .B(n4167), .C(n4168), .D(n4169), .Z(U3_U13_Z_9) );
  AO2 U4658 ( .A(n4160), .B(n4507), .C(n4151), .D(rEIP[9]), .Z(n4169) );
  ND2 U4659 ( .A(n4170), .B(n2195), .Z(n4168) );
  AO3 U4660 ( .A(n4502), .B(n4167), .C(n4171), .D(n4172), .Z(U3_U13_Z_8) );
  AO2 U4661 ( .A(n4160), .B(n4503), .C(n4151), .D(rEIP[8]), .Z(n4172) );
  ND2 U4662 ( .A(n4170), .B(n2196), .Z(n4171) );
  AO3 U4663 ( .A(n4497), .B(n4167), .C(n4173), .D(n4174), .Z(U3_U13_Z_7) );
  AO2 U4664 ( .A(n4160), .B(n4499), .C(n4151), .D(rEIP[7]), .Z(n4174) );
  ND2 U4665 ( .A(n4498), .B(n4170), .Z(n4173) );
  AO3 U4666 ( .A(n4492), .B(n4167), .C(n4175), .D(n4176), .Z(U3_U13_Z_6) );
  AO2 U4667 ( .A(n4160), .B(n4494), .C(n4151), .D(rEIP[6]), .Z(n4176) );
  ND2 U4668 ( .A(n4493), .B(n4170), .Z(n4175) );
  AO3 U4669 ( .A(n4487), .B(n4167), .C(n4177), .D(n4178), .Z(U3_U13_Z_5) );
  AO2 U4670 ( .A(n4160), .B(n4489), .C(n4151), .D(rEIP[5]), .Z(n4178) );
  ND2 U4671 ( .A(n4488), .B(n4170), .Z(n4177) );
  AO3 U4672 ( .A(n4482), .B(n4167), .C(n4179), .D(n4180), .Z(U3_U13_Z_4) );
  AO2 U4673 ( .A(n4160), .B(n4484), .C(n4151), .D(rEIP[4]), .Z(n4180) );
  ND2 U4674 ( .A(n4483), .B(n4170), .Z(n4179) );
  AO3 U4675 ( .A(n4647), .B(n4167), .C(n4181), .D(n4182), .Z(U3_U13_Z_31) );
  AO2 U4676 ( .A(n4160), .B(n2197), .C(n4151), .D(rEIP[31]), .Z(n4182) );
  ND2 U4677 ( .A(n4657), .B(n4170), .Z(n4181) );
  AO3 U4678 ( .A(n4644), .B(n4167), .C(n4183), .D(n4184), .Z(U3_U13_Z_30) );
  AO2 U4679 ( .A(n4160), .B(n2198), .C(n4151), .D(rEIP[30]), .Z(n4184) );
  ND2 U4680 ( .A(n4645), .B(n4170), .Z(n4183) );
  AO3 U4681 ( .A(n4477), .B(n4167), .C(n4185), .D(n4186), .Z(U3_U13_Z_3) );
  AO2 U4682 ( .A(n4160), .B(n4479), .C(n4151), .D(rEIP[3]), .Z(n4186) );
  ND2 U4683 ( .A(n4478), .B(n4170), .Z(n4185) );
  AO3 U4684 ( .A(n4587), .B(n4167), .C(n4187), .D(n4188), .Z(U3_U13_Z_29) );
  AO2 U4685 ( .A(n4160), .B(n2199), .C(n4151), .D(rEIP[29]), .Z(n4188) );
  ND2 U4686 ( .A(n4588), .B(n4170), .Z(n4187) );
  AO3 U4687 ( .A(n4583), .B(n4167), .C(n4189), .D(n4190), .Z(U3_U13_Z_28) );
  AO2 U4688 ( .A(n4160), .B(n2200), .C(n4151), .D(rEIP[28]), .Z(n4190) );
  ND2 U4689 ( .A(n4584), .B(n4170), .Z(n4189) );
  AO3 U4690 ( .A(n4579), .B(n4167), .C(n4191), .D(n4192), .Z(U3_U13_Z_27) );
  AO2 U4691 ( .A(n4160), .B(n2201), .C(n4151), .D(rEIP[27]), .Z(n4192) );
  ND2 U4692 ( .A(n4580), .B(n4170), .Z(n4191) );
  AO3 U4693 ( .A(n4575), .B(n4167), .C(n4193), .D(n4194), .Z(U3_U13_Z_26) );
  AO2 U4694 ( .A(n4160), .B(n2202), .C(n4151), .D(rEIP[26]), .Z(n4194) );
  ND2 U4695 ( .A(n4576), .B(n4170), .Z(n4193) );
  AO3 U4696 ( .A(n4571), .B(n4167), .C(n4195), .D(n4196), .Z(U3_U13_Z_25) );
  AO2 U4697 ( .A(n4160), .B(n2203), .C(n4151), .D(rEIP[25]), .Z(n4196) );
  ND2 U4698 ( .A(n4572), .B(n4170), .Z(n4195) );
  AO3 U4699 ( .A(n4567), .B(n4167), .C(n4197), .D(n4198), .Z(U3_U13_Z_24) );
  AO2 U4700 ( .A(n4160), .B(n2204), .C(n4151), .D(rEIP[24]), .Z(n4198) );
  ND2 U4701 ( .A(n4568), .B(n4170), .Z(n4197) );
  AO3 U4702 ( .A(n4563), .B(n4167), .C(n4199), .D(n4200), .Z(U3_U13_Z_23) );
  AO2 U4703 ( .A(n4160), .B(n2205), .C(n4151), .D(rEIP[23]), .Z(n4200) );
  ND2 U4704 ( .A(n4564), .B(n4170), .Z(n4199) );
  AO3 U4705 ( .A(n4559), .B(n4167), .C(n4201), .D(n4202), .Z(U3_U13_Z_22) );
  AO2 U4706 ( .A(n4160), .B(n4557), .C(n4151), .D(rEIP[22]), .Z(n4202) );
  ND2 U4707 ( .A(n4560), .B(n4170), .Z(n4201) );
  AO3 U4708 ( .A(n4555), .B(n4167), .C(n4203), .D(n4204), .Z(U3_U13_Z_21) );
  AO2 U4709 ( .A(n4160), .B(n4553), .C(n4151), .D(rEIP[21]), .Z(n4204) );
  ND2 U4710 ( .A(n4556), .B(n4170), .Z(n4203) );
  AO3 U4711 ( .A(n4551), .B(n4167), .C(n4205), .D(n4206), .Z(U3_U13_Z_20) );
  AO2 U4712 ( .A(n4160), .B(n4549), .C(n4151), .D(rEIP[20]), .Z(n4206) );
  ND2 U4713 ( .A(n4552), .B(n4170), .Z(n4205) );
  AO3 U4714 ( .A(n4472), .B(n4167), .C(n4207), .D(n4208), .Z(U3_U13_Z_2) );
  AO2 U4715 ( .A(n4160), .B(n4474), .C(n4151), .D(rEIP[2]), .Z(n4208) );
  ND2 U4716 ( .A(n4473), .B(n4170), .Z(n4207) );
  AO3 U4717 ( .A(n4547), .B(n4167), .C(n4209), .D(n4210), .Z(U3_U13_Z_19) );
  AO2 U4718 ( .A(n4160), .B(n4545), .C(n4151), .D(rEIP[19]), .Z(n4210) );
  ND2 U4719 ( .A(n4548), .B(n4170), .Z(n4209) );
  AO3 U4720 ( .A(n4543), .B(n4167), .C(n4211), .D(n4212), .Z(U3_U13_Z_18) );
  AO2 U4721 ( .A(n4160), .B(n4541), .C(n4151), .D(rEIP[18]), .Z(n4212) );
  ND2 U4722 ( .A(n4544), .B(n4170), .Z(n4211) );
  AO3 U4723 ( .A(n4539), .B(n4167), .C(n4213), .D(n4214), .Z(U3_U13_Z_17) );
  AO2 U4724 ( .A(n4160), .B(n4537), .C(n4151), .D(rEIP[17]), .Z(n4214) );
  ND2 U4725 ( .A(n4540), .B(n4170), .Z(n4213) );
  AO3 U4726 ( .A(n4535), .B(n4167), .C(n4215), .D(n4216), .Z(U3_U13_Z_16) );
  AO2 U4727 ( .A(n4160), .B(n4533), .C(n4151), .D(rEIP[16]), .Z(n4216) );
  ND2 U4728 ( .A(n4536), .B(n4170), .Z(n4215) );
  AO3 U4729 ( .A(n4530), .B(n4167), .C(n4217), .D(n4218), .Z(U3_U13_Z_15) );
  AO2 U4730 ( .A(n4160), .B(n4531), .C(n4151), .D(rEIP[15]), .Z(n4218) );
  ND2 U4731 ( .A(n4170), .B(n2206), .Z(n4217) );
  AO3 U4732 ( .A(n4526), .B(n4167), .C(n4219), .D(n4220), .Z(U3_U13_Z_14) );
  AO2 U4733 ( .A(n4160), .B(n4527), .C(n4151), .D(rEIP[14]), .Z(n4220) );
  ND2 U4734 ( .A(n4170), .B(n2207), .Z(n4219) );
  AO3 U4735 ( .A(n4522), .B(n4167), .C(n4221), .D(n4222), .Z(U3_U13_Z_13) );
  AO2 U4736 ( .A(n4160), .B(n4523), .C(n4151), .D(rEIP[13]), .Z(n4222) );
  ND2 U4737 ( .A(n4170), .B(n2208), .Z(n4221) );
  AO3 U4738 ( .A(n4518), .B(n4167), .C(n4223), .D(n4224), .Z(U3_U13_Z_12) );
  AO2 U4739 ( .A(n4160), .B(n4519), .C(n4151), .D(rEIP[12]), .Z(n4224) );
  ND2 U4740 ( .A(n4170), .B(n2209), .Z(n4223) );
  AO3 U4741 ( .A(n4514), .B(n4167), .C(n4225), .D(n4226), .Z(U3_U13_Z_11) );
  AO2 U4742 ( .A(n4160), .B(n4515), .C(n4151), .D(rEIP[11]), .Z(n4226) );
  ND2 U4743 ( .A(n4170), .B(n2210), .Z(n4225) );
  AO3 U4744 ( .A(n4510), .B(n4167), .C(n4227), .D(n4228), .Z(U3_U13_Z_10) );
  AO2 U4745 ( .A(n4160), .B(n4511), .C(n4151), .D(rEIP[10]), .Z(n4228) );
  ND2 U4746 ( .A(n4170), .B(n2211), .Z(n4227) );
  AO3 U4747 ( .A(n4459), .B(n4167), .C(n4229), .D(n4230), .Z(U3_U13_Z_1) );
  AO2 U4748 ( .A(n4160), .B(n4469), .C(n4151), .D(rEIP[1]), .Z(n4230) );
  ND2 U4749 ( .A(n4453), .B(n4170), .Z(n4229) );
  AO3 U4750 ( .A(n4460), .B(n4167), .C(n4231), .D(n4232), .Z(U3_U13_Z_0) );
  AO2 U4751 ( .A(n4160), .B(n4465), .C(n4151), .D(rEIP[0]), .Z(n4232) );
  NR3 U4752 ( .A(n2214), .B(n2359), .C(n3582), .Z(n4151) );
  ND3 U4753 ( .A(n3805), .B(n2286), .C(n2552), .Z(n3582) );
  IV U4754 ( .A(n2395), .Z(n2552) );
  NR2 U4755 ( .A(n2776), .B(n2359), .Z(n4160) );
  ND2 U4756 ( .A(n4006), .B(n4033), .Z(n2776) );
  AN3 U4757 ( .A(n3541), .B(n3556), .C(n4035), .Z(n4006) );
  NR4 U4758 ( .A(n3564), .B(n4233), .C(n4234), .D(n4235), .Z(n4035) );
  ND2 U4759 ( .A(n4654), .B(n4170), .Z(n4231) );
  ND3 U4760 ( .A(n4010), .B(n4143), .C(n4153), .Z(n4170) );
  AO6 U4761 ( .A(n2286), .B(n3870), .C(n4030), .Z(n4153) );
  NR2 U4762 ( .A(n3805), .B(n3587), .Z(n4030) );
  IV U4763 ( .A(n3795), .Z(n3870) );
  ND2 U4764 ( .A(n3864), .B(n2284), .Z(n3795) );
  IV U4765 ( .A(n2287), .Z(n2284) );
  NR2 U4766 ( .A(n2315), .B(n2309), .Z(n2287) );
  NR3 U4767 ( .A(n4666), .B(n4651), .C(n2150), .Z(n2309) );
  AN3 U4768 ( .A(n2150), .B(n2212), .C(n4651), .Z(n2315) );
  IV U4769 ( .A(n3583), .Z(n3864) );
  ND2 U4770 ( .A(n2288), .B(n3796), .Z(n3583) );
  IV U4771 ( .A(n2245), .Z(n3796) );
  ND2 U4772 ( .A(n2278), .B(n3805), .Z(n2245) );
  IV U4773 ( .A(n2549), .Z(n2288) );
  IV U4774 ( .A(READY_n), .Z(n2286) );
  AO6 U4775 ( .A(n2278), .B(n3810), .C(n3826), .Z(n4143) );
  IV U4776 ( .A(n3812), .Z(n3826) );
  ND2 U4777 ( .A(n2278), .B(n2613), .Z(n3812) );
  IV U4778 ( .A(n2615), .Z(n2613) );
  NR2 U4779 ( .A(n2254), .B(n4031), .Z(n2615) );
  NR2 U4780 ( .A(n2772), .B(n2371), .Z(n4031) );
  IV U4781 ( .A(n4008), .Z(n2254) );
  ND2 U4782 ( .A(n3685), .B(n3805), .Z(n4008) );
  IV U4783 ( .A(n2371), .Z(n3805) );
  IV U4784 ( .A(n2724), .Z(n3685) );
  NR2 U4785 ( .A(n4236), .B(n2371), .Z(n3810) );
  IV U4786 ( .A(n2359), .Z(n2278) );
  IV U4787 ( .A(U3_U14_Z_7), .Z(n4010) );
  NR2 U4788 ( .A(n3587), .B(n2371), .Z(U3_U14_Z_7) );
  MUX21L U4789 ( .A(n3683), .B(n4237), .S(n4238), .Z(n2371) );
  AO2 U4790 ( .A(n3809), .B(n4011), .C(n4239), .D(n2372), .Z(n4238) );
  AO1 U4791 ( .A(n3940), .B(n2578), .C(n4240), .D(n4241), .Z(n4011) );
  MUX21L U4792 ( .A(n4242), .B(n4243), .S(n2167), .Z(n4241) );
  NR2 U4793 ( .A(n4005), .B(n4077), .Z(n4240) );
  AO7 U4794 ( .A(n4632), .B(n2347), .C(n4244), .Z(n3940) );
  IV U4795 ( .A(n4245), .Z(n4244) );
  AO4 U4796 ( .A(n3943), .B(n4382), .C(n2349), .D(n4383), .Z(n4245) );
  AO1 U4797 ( .A(n4246), .B(n4247), .C(n3683), .D(n4248), .Z(n4237) );
  NR3 U4798 ( .A(n4249), .B(n3804), .C(n4250), .Z(n4248) );
  AO2 U4799 ( .A(n2244), .B(n4251), .C(n3804), .D(n4250), .Z(n4247) );
  AO7 U4800 ( .A(n4454), .B(n2145), .C(n4252), .Z(n4251) );
  NR2 U4801 ( .A(n4249), .B(n4253), .Z(n4246) );
  IV U4802 ( .A(n2372), .Z(n3683) );
  ND2 U4803 ( .A(n3804), .B(n2244), .Z(n2372) );
  AN3 U4804 ( .A(n2549), .B(n2395), .C(n2429), .Z(n2244) );
  IV U4805 ( .A(n3684), .Z(n2429) );
  ND2 U4806 ( .A(n3808), .B(n2283), .Z(n3684) );
  ND3 U4807 ( .A(n4254), .B(n3544), .C(n4255), .Z(n2283) );
  ND2 U4808 ( .A(n4033), .B(n4255), .Z(n3808) );
  AN3 U4809 ( .A(n4256), .B(n3553), .C(n4234), .Z(n4255) );
  IV U4810 ( .A(n3550), .Z(n4234) );
  ND2 U4811 ( .A(n4007), .B(n4257), .Z(n2395) );
  ND3 U4812 ( .A(n4258), .B(n3547), .C(n4257), .Z(n2549) );
  NR3 U4813 ( .A(n4233), .B(n4259), .C(n4260), .Z(n4257) );
  IV U4814 ( .A(n3559), .Z(n4233) );
  AN3 U4815 ( .A(n2772), .B(n2724), .C(n4236), .Z(n3804) );
  IV U4816 ( .A(n3682), .Z(n4236) );
  NR2 U4817 ( .A(n4261), .B(n4254), .Z(n3682) );
  ND2 U4818 ( .A(n4262), .B(n4007), .Z(n2724) );
  NR2 U4819 ( .A(n3547), .B(n3544), .Z(n4007) );
  ND2 U4820 ( .A(n4262), .B(n4033), .Z(n2772) );
  NR2 U4821 ( .A(n4254), .B(n4258), .Z(n4033) );
  IV U4822 ( .A(n3547), .Z(n4254) );
  NR3 U4823 ( .A(n3559), .B(n4260), .C(n3556), .Z(n4262) );
  ND4 U4824 ( .A(n4235), .B(n4034), .C(n3564), .D(n3550), .Z(n4260) );
  IV U4825 ( .A(n3541), .Z(n4034) );
  IV U4826 ( .A(n3809), .Z(n3587) );
  NR4 U4827 ( .A(n2359), .B(n2387), .C(n4263), .D(n4239), .Z(n3809) );
  AO2 U4828 ( .A(n4467), .B(n4264), .C(n2171), .D(n4265), .Z(n4239) );
  OR2 U4829 ( .A(n4264), .B(n4467), .Z(n4265) );
  AO1 U4830 ( .A(n4253), .B(n4266), .C(n4249), .D(n4250), .Z(n4263) );
  EO U4831 ( .A(n4267), .B(n4268), .Z(n4250) );
  EO U4832 ( .A(n4456), .B(n4653), .Z(n4267) );
  EO U4833 ( .A(n4264), .B(n4269), .Z(n4249) );
  ND2 U4834 ( .A(n4467), .B(n2171), .Z(n4269) );
  AO2 U4835 ( .A(n2148), .B(n4268), .C(n4270), .D(n4456), .Z(n4264) );
  OR2 U4836 ( .A(n4268), .B(n2148), .Z(n4270) );
  AO2 U4837 ( .A(n4252), .B(n4461), .C(n2146), .D(n4271), .Z(n4268) );
  OR2 U4838 ( .A(n4461), .B(n4252), .Z(n4271) );
  EO U4839 ( .A(n2145), .B(n2169), .Z(n4266) );
  EN U4840 ( .A(n4272), .B(n4252), .Z(n4253) );
  ND2 U4841 ( .A(n4454), .B(n2145), .Z(n4252) );
  EO U4842 ( .A(n4455), .B(n4461), .Z(n4272) );
  IV U4843 ( .A(n3586), .Z(n2387) );
  NR2 U4844 ( .A(n4261), .B(n3547), .Z(n3586) );
  AO3 U4845 ( .A(n4156), .B(n2570), .C(n4273), .D(n4274), .Z(n3547) );
  AO2 U4846 ( .A(n2571), .B(n4159), .C(n2578), .D(n3834), .Z(n4274) );
  OR2 U4847 ( .A(n4275), .B(n4276), .Z(n3834) );
  AO4 U4848 ( .A(n4277), .B(n4421), .C(n3943), .D(n4422), .Z(n4276) );
  AO4 U4849 ( .A(n2349), .B(n4423), .C(n2347), .D(n4597), .Z(n4275) );
  OR2 U4850 ( .A(n4278), .B(n4279), .Z(n4159) );
  AO4 U4851 ( .A(n4277), .B(n4427), .C(n3943), .D(n4428), .Z(n4279) );
  AO4 U4852 ( .A(n2349), .B(n4429), .C(n2347), .D(n4599), .Z(n4278) );
  AO7 U4853 ( .A(n4280), .B(n4281), .C(n3820), .Z(n4273) );
  AO4 U4854 ( .A(n4424), .B(n2347), .C(n4596), .D(n2349), .Z(n4281) );
  AO4 U4855 ( .A(n4425), .B(n3943), .C(n4426), .D(n4277), .Z(n4280) );
  NR2 U4856 ( .A(n4282), .B(n4283), .Z(n4156) );
  AO4 U4857 ( .A(n4277), .B(n4418), .C(n3943), .D(n4419), .Z(n4283) );
  AO4 U4858 ( .A(n2349), .B(n4420), .C(n2347), .D(n4598), .Z(n4282) );
  ND4 U4859 ( .A(n4256), .B(n4235), .C(n4258), .D(n3550), .Z(n4261) );
  AO3 U4860 ( .A(n4146), .B(n2570), .C(n4284), .D(n4285), .Z(n3550) );
  AO2 U4861 ( .A(n2571), .B(n4149), .C(n2578), .D(n3828), .Z(n4285) );
  OR2 U4862 ( .A(n4286), .B(n4287), .Z(n3828) );
  AO4 U4863 ( .A(n4277), .B(n4399), .C(n3943), .D(n4400), .Z(n4287) );
  AO4 U4864 ( .A(n2349), .B(n4401), .C(n2347), .D(n4603), .Z(n4286) );
  OR2 U4865 ( .A(n4288), .B(n4289), .Z(n4149) );
  AO4 U4866 ( .A(n4277), .B(n4404), .C(n3943), .D(n4405), .Z(n4289) );
  AO4 U4867 ( .A(n2349), .B(n4601), .C(n2347), .D(n4605), .Z(n4288) );
  AO7 U4868 ( .A(n4290), .B(n4291), .C(n3820), .Z(n4284) );
  AO4 U4869 ( .A(n4402), .B(n2347), .C(n4602), .D(n2349), .Z(n4291) );
  AO4 U4870 ( .A(n4664), .B(n3943), .C(n4403), .D(n4277), .Z(n4290) );
  NR2 U4871 ( .A(n4292), .B(n4293), .Z(n4146) );
  AO4 U4872 ( .A(n4277), .B(n4396), .C(n3943), .D(n4397), .Z(n4293) );
  AO4 U4873 ( .A(n2349), .B(n4398), .C(n2347), .D(n4604), .Z(n4292) );
  IV U4874 ( .A(n3544), .Z(n4258) );
  AO3 U4875 ( .A(n4163), .B(n2570), .C(n4294), .D(n4295), .Z(n3544) );
  AO2 U4876 ( .A(n2571), .B(n4166), .C(n2578), .D(n3841), .Z(n4295) );
  OR2 U4877 ( .A(n4296), .B(n4297), .Z(n3841) );
  AO4 U4878 ( .A(n4277), .B(n4409), .C(n3943), .D(n4410), .Z(n4297) );
  AO4 U4879 ( .A(n2349), .B(n4411), .C(n2347), .D(n4592), .Z(n4296) );
  OR2 U4880 ( .A(n4298), .B(n4299), .Z(n4166) );
  AO4 U4881 ( .A(n4277), .B(n4415), .C(n3943), .D(n4416), .Z(n4299) );
  AO4 U4882 ( .A(n2349), .B(n4417), .C(n2347), .D(n4594), .Z(n4298) );
  AO7 U4883 ( .A(n4300), .B(n4301), .C(n3820), .Z(n4294) );
  AO4 U4884 ( .A(n4412), .B(n2347), .C(n4591), .D(n2349), .Z(n4301) );
  AO4 U4885 ( .A(n4413), .B(n3943), .C(n4414), .D(n4277), .Z(n4300) );
  NR2 U4886 ( .A(n4302), .B(n4303), .Z(n4163) );
  AO4 U4887 ( .A(n4277), .B(n4406), .C(n3943), .D(n4407), .Z(n4303) );
  AO4 U4888 ( .A(n2349), .B(n4408), .C(n2347), .D(n4593), .Z(n4302) );
  IV U4889 ( .A(n3553), .Z(n4235) );
  AO3 U4890 ( .A(n4141), .B(n2570), .C(n4304), .D(n4305), .Z(n3553) );
  AO2 U4891 ( .A(n2571), .B(n4140), .C(n2578), .D(n4108), .Z(n4305) );
  IV U4892 ( .A(n3819), .Z(n4108) );
  NR2 U4893 ( .A(n4306), .B(n4307), .Z(n3819) );
  AO4 U4894 ( .A(n4277), .B(n4432), .C(n3943), .D(n4433), .Z(n4307) );
  AO4 U4895 ( .A(n2349), .B(n4434), .C(n2347), .D(n4609), .Z(n4306) );
  OR2 U4896 ( .A(n4308), .B(n4309), .Z(n4140) );
  AO4 U4897 ( .A(n4277), .B(n4437), .C(n3943), .D(n4438), .Z(n4309) );
  AO4 U4898 ( .A(n2349), .B(n4439), .C(n2347), .D(n4611), .Z(n4308) );
  AO7 U4899 ( .A(n4310), .B(n4311), .C(n3820), .Z(n4304) );
  AO4 U4900 ( .A(n4435), .B(n2347), .C(n4608), .D(n2349), .Z(n4311) );
  AO4 U4901 ( .A(n4663), .B(n3943), .C(n4436), .D(n4277), .Z(n4310) );
  NR2 U4902 ( .A(n4312), .B(n4313), .Z(n4141) );
  AO4 U4903 ( .A(n4277), .B(n4430), .C(n3943), .D(n4431), .Z(n4313) );
  AO4 U4904 ( .A(n2349), .B(n4607), .C(n2347), .D(n4610), .Z(n4312) );
  NR4 U4905 ( .A(n3564), .B(n3559), .C(n3541), .D(n4259), .Z(n4256) );
  IV U4906 ( .A(n3556), .Z(n4259) );
  AO3 U4907 ( .A(n4136), .B(n2570), .C(n4314), .D(n4315), .Z(n3556) );
  AO2 U4908 ( .A(n2571), .B(n4135), .C(n2578), .D(n4100), .Z(n4315) );
  IV U4909 ( .A(n3909), .Z(n4100) );
  NR2 U4910 ( .A(n4316), .B(n4317), .Z(n3909) );
  AO4 U4911 ( .A(n4277), .B(n4442), .C(n3943), .D(n4443), .Z(n4317) );
  AO4 U4912 ( .A(n2349), .B(n4444), .C(n2347), .D(n4615), .Z(n4316) );
  OR2 U4913 ( .A(n4318), .B(n4319), .Z(n4135) );
  AO4 U4914 ( .A(n4277), .B(n4447), .C(n3943), .D(n4448), .Z(n4319) );
  AO4 U4915 ( .A(n2349), .B(n4449), .C(n2347), .D(n4617), .Z(n4318) );
  AO7 U4916 ( .A(n4320), .B(n4321), .C(n3820), .Z(n4314) );
  AO4 U4917 ( .A(n4445), .B(n2347), .C(n4614), .D(n2349), .Z(n4321) );
  AO4 U4918 ( .A(n4662), .B(n3943), .C(n4446), .D(n4277), .Z(n4320) );
  NR2 U4919 ( .A(n4322), .B(n4323), .Z(n4136) );
  AO4 U4920 ( .A(n4277), .B(n4440), .C(n3943), .D(n4441), .Z(n4323) );
  AO4 U4921 ( .A(n2349), .B(n4613), .C(n2347), .D(n4616), .Z(n4322) );
  AO3 U4922 ( .A(n4077), .B(n2570), .C(n4324), .D(n4325), .Z(n3541) );
  EO1 U4923 ( .A(n2578), .B(n3885), .C(n4005), .D(n4242), .Z(n4325) );
  NR2 U4924 ( .A(n4326), .B(n4327), .Z(n4242) );
  AO4 U4925 ( .A(n4277), .B(n4384), .C(n3943), .D(n4385), .Z(n4327) );
  AO4 U4926 ( .A(n2349), .B(n4386), .C(n2347), .D(n4635), .Z(n4326) );
  IV U4927 ( .A(n4243), .Z(n3885) );
  NR2 U4928 ( .A(n4328), .B(n4329), .Z(n4243) );
  AO4 U4929 ( .A(n4277), .B(n4379), .C(n3943), .D(n4380), .Z(n4329) );
  AO4 U4930 ( .A(n2349), .B(n4381), .C(n2347), .D(n4633), .Z(n4328) );
  AO7 U4931 ( .A(n4330), .B(n4331), .C(n3820), .Z(n4324) );
  AO4 U4932 ( .A(n4382), .B(n2347), .C(n4632), .D(n2349), .Z(n4331) );
  AO4 U4933 ( .A(n4659), .B(n3943), .C(n4383), .D(n4277), .Z(n4330) );
  NR2 U4934 ( .A(n4332), .B(n4333), .Z(n4077) );
  AO4 U4935 ( .A(n4277), .B(n4376), .C(n3943), .D(n4377), .Z(n4333) );
  AO4 U4936 ( .A(n2349), .B(n4378), .C(n2347), .D(n4634), .Z(n4332) );
  AO3 U4937 ( .A(n4131), .B(n2570), .C(n4334), .D(n4335), .Z(n3559) );
  AO2 U4938 ( .A(n2571), .B(n4130), .C(n2578), .D(n4092), .Z(n4335) );
  IV U4939 ( .A(n3901), .Z(n4092) );
  NR2 U4940 ( .A(n4336), .B(n4337), .Z(n3901) );
  AO4 U4941 ( .A(n4277), .B(n4368), .C(n3943), .D(n4369), .Z(n4337) );
  AO4 U4942 ( .A(n2349), .B(n4370), .C(n2347), .D(n4621), .Z(n4336) );
  OR2 U4943 ( .A(n4338), .B(n4339), .Z(n4130) );
  AO4 U4944 ( .A(n4277), .B(n4373), .C(n3943), .D(n4374), .Z(n4339) );
  AO4 U4945 ( .A(n2349), .B(n4375), .C(n2347), .D(n4623), .Z(n4338) );
  AO7 U4946 ( .A(n4340), .B(n4341), .C(n3820), .Z(n4334) );
  AO4 U4947 ( .A(n4371), .B(n2347), .C(n4620), .D(n2349), .Z(n4341) );
  AO4 U4948 ( .A(n4661), .B(n3943), .C(n4372), .D(n4277), .Z(n4340) );
  NR2 U4949 ( .A(n4342), .B(n4343), .Z(n4131) );
  AO4 U4950 ( .A(n4277), .B(n4366), .C(n3943), .D(n4367), .Z(n4343) );
  AO4 U4951 ( .A(n2349), .B(n4619), .C(n2347), .D(n4622), .Z(n4342) );
  AO3 U4952 ( .A(n4126), .B(n2570), .C(n4344), .D(n4345), .Z(n3564) );
  AO2 U4953 ( .A(n2571), .B(n4125), .C(n2578), .D(n4084), .Z(n4345) );
  IV U4954 ( .A(n3893), .Z(n4084) );
  NR2 U4955 ( .A(n4346), .B(n4347), .Z(n3893) );
  AO4 U4956 ( .A(n4277), .B(n4389), .C(n3943), .D(n4390), .Z(n4347) );
  AO4 U4957 ( .A(n2349), .B(n4391), .C(n2347), .D(n4628), .Z(n4346) );
  IV U4958 ( .A(n2348), .Z(n2578) );
  ND2 U4959 ( .A(n2167), .B(n2145), .Z(n2348) );
  OR2 U4960 ( .A(n4348), .B(n4349), .Z(n4125) );
  AO4 U4961 ( .A(n4277), .B(n4394), .C(n3943), .D(n4395), .Z(n4349) );
  AO4 U4962 ( .A(n2349), .B(n4626), .C(n2347), .D(n4630), .Z(n4348) );
  IV U4963 ( .A(n4005), .Z(n2571) );
  ND2 U4964 ( .A(n4461), .B(n2145), .Z(n4005) );
  AO7 U4965 ( .A(n4350), .B(n4351), .C(n3820), .Z(n4344) );
  IV U4966 ( .A(n2610), .Z(n3820) );
  ND2 U4967 ( .A(n4461), .B(n4468), .Z(n2610) );
  AO4 U4968 ( .A(n4392), .B(n2347), .C(n4627), .D(n2349), .Z(n4351) );
  AO4 U4969 ( .A(n4660), .B(n3943), .C(n4393), .D(n4277), .Z(n4350) );
  ND2 U4970 ( .A(n4468), .B(n2167), .Z(n2570) );
  NR2 U4971 ( .A(n4352), .B(n4353), .Z(n4126) );
  AO4 U4972 ( .A(n4277), .B(n4387), .C(n3943), .D(n4388), .Z(n4353) );
  ND2 U4973 ( .A(n4467), .B(n4653), .Z(n3943) );
  ND2 U4974 ( .A(n2148), .B(n2213), .Z(n4277) );
  AO4 U4975 ( .A(n2349), .B(n4625), .C(n2347), .D(n4629), .Z(n4352) );
  ND2 U4976 ( .A(n4467), .B(n2148), .Z(n2347) );
  ND2 U4977 ( .A(n4653), .B(n2213), .Z(n2349) );
  OR3 U4978 ( .A(n4450), .B(n4658), .C(n2396), .Z(n2359) );
  AN2 U4979 ( .A(n3540), .B(n2590), .Z(n4167) );
  ND2 U4980 ( .A(n2618), .B(n2214), .Z(n2590) );
  NR2 U4981 ( .A(n2389), .B(n2617), .Z(n3540) );
  IV U4982 ( .A(n2360), .Z(n2617) );
  OR3 U4983 ( .A(n4450), .B(n2396), .C(n2151), .Z(n2360) );
  ND2 U4984 ( .A(n4458), .B(n4668), .Z(n2396) );
  IV U4985 ( .A(n2598), .Z(n2389) );
  ND2 U4986 ( .A(n2618), .B(n4665), .Z(n2598) );
  IV U4987 ( .A(n2556), .Z(n2618) );
  ND2 U4988 ( .A(n2390), .B(n3565), .Z(n2556) );
  IV U4989 ( .A(n3760), .Z(n3565) );
  ND2 U4990 ( .A(n4658), .B(n4450), .Z(n3760) );
  NR2 U4991 ( .A(n2183), .B(n4668), .Z(n2390) );
  EO r1165_U53 ( .A(n2140), .B(U3_U7_Z_0), .Z(N2787) );
  AN2 r1165_U52 ( .A(n2140), .B(U3_U7_Z_0), .Z(r1165_n15) );
  EO r1165_U51 ( .A(U3_U8_Z_1), .B(U3_U7_Z_1), .Z(r1165_n17) );
  EO r1165_U50 ( .A(r1165_n15), .B(r1165_n17), .Z(N2788) );
  OR2 r1165_U49 ( .A(r1165_n15), .B(U3_U7_Z_1), .Z(r1165_n16) );
  AO2 r1165_U48 ( .A(r1165_n15), .B(U3_U7_Z_1), .C(r1165_n16), .D(U3_U8_Z_1), 
        .Z(r1165_n13) );
  EN r1165_U47 ( .A(U3_U8_Z_2), .B(U3_U7_Z_2), .Z(r1165_n14) );
  EO r1165_U46 ( .A(r1165_n13), .B(r1165_n14), .Z(N2789) );
  IV r1165_U45 ( .A(r1165_n13), .Z(r1165_n11) );
  OR2 r1165_U44 ( .A(U3_U7_Z_2), .B(r1165_n11), .Z(r1165_n12) );
  AO2 r1165_U43 ( .A(r1165_n11), .B(U3_U7_Z_2), .C(r1165_n12), .D(U3_U8_Z_2), 
        .Z(r1165_n9) );
  EN r1165_U42 ( .A(U3_U8_Z_3), .B(U3_U7_Z_3), .Z(r1165_n10) );
  EO r1165_U41 ( .A(r1165_n9), .B(r1165_n10), .Z(N2790) );
  IV r1165_U40 ( .A(r1165_n9), .Z(r1165_n7) );
  AN2 r1165_U39 ( .A(r1165_n7), .B(U3_U7_Z_3), .Z(r1165_n8) );
  AO4 r1165_U38 ( .A(U3_U7_Z_3), .B(r1165_n7), .C(U3_U8_Z_3), .D(r1165_n8), 
        .Z(r1165_n6) );
  IV r1165_U37 ( .A(U3_U8_Z_4), .Z(r1165_n5) );
  EO r1165_U36 ( .A(r1165_n6), .B(r1165_n5), .Z(N2791) );
  NR2 r1165_U35 ( .A(r1165_n5), .B(r1165_n6), .Z(r1165_n4) );
  EO r1165_U34 ( .A(U3_U8_Z_5), .B(r1165_n4), .Z(N2792) );
  ND2 r1165_U33 ( .A(U3_U8_Z_5), .B(r1165_n4), .Z(r1165_n2) );
  IV r1165_U32 ( .A(U3_U8_Z_6), .Z(r1165_n3) );
  EO r1165_U31 ( .A(r1165_n2), .B(r1165_n3), .Z(N818) );
  NR2 r1165_U30 ( .A(r1165_n2), .B(r1165_n3), .Z(r1165_n1) );
  EO r1165_U29 ( .A(U3_U8_Z_7), .B(r1165_n1), .Z(N819) );
  EO r1164_U352 ( .A(U3_U6_Z_0), .B(U3_U5_Z_0), .Z(N2579) );
  EN r1164_U351 ( .A(U3_U6_Z_10), .B(U3_U5_Z_10), .Z(r1164_n129) );
  AN2 r1164_U350 ( .A(U3_U5_Z_0), .B(U3_U6_Z_0), .Z(r1164_n145) );
  AO5 r1164_U349 ( .A(U3_U5_Z_1), .B(U3_U6_Z_1), .C(r1164_n145), .Z(r1164_n27)
         );
  IV r1164_U348 ( .A(r1164_n27), .Z(r1164_n143) );
  OR2 r1164_U347 ( .A(r1164_n143), .B(U3_U5_Z_2), .Z(r1164_n144) );
  AO2 r1164_U346 ( .A(r1164_n143), .B(U3_U5_Z_2), .C(r1164_n144), .D(U3_U6_Z_2), .Z(r1164_n16) );
  IV r1164_U345 ( .A(r1164_n16), .Z(r1164_n141) );
  OR2 r1164_U344 ( .A(U3_U5_Z_3), .B(r1164_n141), .Z(r1164_n142) );
  AO2 r1164_U343 ( .A(r1164_n141), .B(U3_U5_Z_3), .C(r1164_n142), .D(U3_U6_Z_3), .Z(r1164_n14) );
  IV r1164_U342 ( .A(r1164_n14), .Z(r1164_n139) );
  AN2 r1164_U341 ( .A(r1164_n139), .B(U3_U5_Z_4), .Z(r1164_n140) );
  AO4 r1164_U340 ( .A(U3_U5_Z_4), .B(r1164_n139), .C(U3_U6_Z_4), .D(r1164_n140), .Z(r1164_n13) );
  IV r1164_U339 ( .A(r1164_n13), .Z(r1164_n137) );
  OR2 r1164_U338 ( .A(r1164_n137), .B(U3_U5_Z_5), .Z(r1164_n138) );
  AO2 r1164_U337 ( .A(r1164_n137), .B(U3_U5_Z_5), .C(r1164_n138), .D(U3_U6_Z_5), .Z(r1164_n10) );
  IV r1164_U336 ( .A(r1164_n10), .Z(r1164_n135) );
  AN2 r1164_U335 ( .A(r1164_n135), .B(U3_U5_Z_6), .Z(r1164_n136) );
  AO4 r1164_U334 ( .A(U3_U5_Z_6), .B(r1164_n135), .C(U3_U6_Z_6), .D(r1164_n136), .Z(r1164_n9) );
  IV r1164_U333 ( .A(r1164_n9), .Z(r1164_n133) );
  OR2 r1164_U332 ( .A(r1164_n133), .B(U3_U5_Z_7), .Z(r1164_n134) );
  AO2 r1164_U331 ( .A(r1164_n133), .B(U3_U5_Z_7), .C(r1164_n134), .D(U3_U6_Z_7), .Z(r1164_n5) );
  IV r1164_U330 ( .A(r1164_n5), .Z(r1164_n3) );
  ND2 r1164_U329 ( .A(U3_U5_Z_8), .B(r1164_n3), .Z(r1164_n131) );
  IV r1164_U328 ( .A(U3_U6_Z_8), .Z(r1164_n132) );
  IV r1164_U327 ( .A(U3_U5_Z_8), .Z(r1164_n6) );
  AO2 r1164_U326 ( .A(r1164_n131), .B(r1164_n132), .C(r1164_n5), .D(r1164_n6), 
        .Z(r1164_n130) );
  AO5 r1164_U325 ( .A(U3_U5_Z_9), .B(U3_U6_Z_9), .C(r1164_n130), .Z(r1164_n128) );
  EO r1164_U324 ( .A(r1164_n129), .B(r1164_n128), .Z(N2589) );
  IV r1164_U323 ( .A(r1164_n128), .Z(r1164_n126) );
  OR2 r1164_U322 ( .A(r1164_n126), .B(U3_U5_Z_10), .Z(r1164_n127) );
  AO2 r1164_U321 ( .A(r1164_n126), .B(U3_U5_Z_10), .C(r1164_n127), .D(
        U3_U6_Z_10), .Z(r1164_n124) );
  EN r1164_U320 ( .A(U3_U6_Z_11), .B(U3_U5_Z_11), .Z(r1164_n125) );
  EO r1164_U319 ( .A(r1164_n124), .B(r1164_n125), .Z(N2590) );
  EN r1164_U318 ( .A(U3_U6_Z_12), .B(U3_U5_Z_12), .Z(r1164_n121) );
  IV r1164_U317 ( .A(r1164_n124), .Z(r1164_n122) );
  AN2 r1164_U316 ( .A(r1164_n122), .B(U3_U5_Z_11), .Z(r1164_n123) );
  AO4 r1164_U315 ( .A(U3_U5_Z_11), .B(r1164_n122), .C(U3_U6_Z_11), .D(
        r1164_n123), .Z(r1164_n120) );
  EO r1164_U314 ( .A(r1164_n121), .B(r1164_n120), .Z(N2591) );
  IV r1164_U313 ( .A(r1164_n120), .Z(r1164_n118) );
  OR2 r1164_U312 ( .A(r1164_n118), .B(U3_U5_Z_12), .Z(r1164_n119) );
  AO2 r1164_U311 ( .A(r1164_n118), .B(U3_U5_Z_12), .C(r1164_n119), .D(
        U3_U6_Z_12), .Z(r1164_n116) );
  EN r1164_U310 ( .A(U3_U6_Z_13), .B(U3_U5_Z_13), .Z(r1164_n117) );
  EO r1164_U309 ( .A(r1164_n116), .B(r1164_n117), .Z(N2592) );
  EN r1164_U308 ( .A(U3_U6_Z_14), .B(U3_U5_Z_14), .Z(r1164_n113) );
  IV r1164_U307 ( .A(r1164_n116), .Z(r1164_n114) );
  AN2 r1164_U306 ( .A(r1164_n114), .B(U3_U5_Z_13), .Z(r1164_n115) );
  AO4 r1164_U305 ( .A(U3_U5_Z_13), .B(r1164_n114), .C(U3_U6_Z_13), .D(
        r1164_n115), .Z(r1164_n112) );
  EO r1164_U304 ( .A(r1164_n113), .B(r1164_n112), .Z(N2593) );
  IV r1164_U303 ( .A(r1164_n112), .Z(r1164_n110) );
  OR2 r1164_U302 ( .A(r1164_n110), .B(U3_U5_Z_14), .Z(r1164_n111) );
  AO2 r1164_U301 ( .A(r1164_n110), .B(U3_U5_Z_14), .C(r1164_n111), .D(
        U3_U6_Z_14), .Z(r1164_n108) );
  EN r1164_U300 ( .A(U3_U6_Z_15), .B(U3_U5_Z_15), .Z(r1164_n109) );
  EO r1164_U299 ( .A(r1164_n108), .B(r1164_n109), .Z(N2594) );
  EN r1164_U298 ( .A(U3_U6_Z_16), .B(U3_U5_Z_16), .Z(r1164_n105) );
  IV r1164_U297 ( .A(r1164_n108), .Z(r1164_n106) );
  AN2 r1164_U296 ( .A(r1164_n106), .B(U3_U5_Z_15), .Z(r1164_n107) );
  AO4 r1164_U295 ( .A(U3_U5_Z_15), .B(r1164_n106), .C(U3_U6_Z_15), .D(
        r1164_n107), .Z(r1164_n104) );
  EO r1164_U294 ( .A(r1164_n105), .B(r1164_n104), .Z(N2595) );
  IV r1164_U293 ( .A(r1164_n104), .Z(r1164_n102) );
  OR2 r1164_U292 ( .A(r1164_n102), .B(U3_U5_Z_16), .Z(r1164_n103) );
  AO2 r1164_U291 ( .A(r1164_n102), .B(U3_U5_Z_16), .C(r1164_n103), .D(
        U3_U6_Z_16), .Z(r1164_n94) );
  IV r1164_U290 ( .A(U3_U6_Z_17), .Z(r1164_n97) );
  EO r1164_U289 ( .A(U3_U5_Z_17), .B(r1164_n97), .Z(r1164_n101) );
  EO r1164_U288 ( .A(r1164_n94), .B(r1164_n101), .Z(N2596) );
  IV r1164_U287 ( .A(U3_U5_Z_18), .Z(r1164_n88) );
  EO r1164_U286 ( .A(r1164_n88), .B(U3_U6_Z_18), .Z(r1164_n99) );
  IV r1164_U285 ( .A(r1164_n94), .Z(r1164_n98) );
  IV r1164_U284 ( .A(U3_U5_Z_17), .Z(r1164_n95) );
  NR2 r1164_U283 ( .A(r1164_n94), .B(r1164_n95), .Z(r1164_n100) );
  AO4 r1164_U282 ( .A(U3_U5_Z_17), .B(r1164_n98), .C(U3_U6_Z_17), .D(
        r1164_n100), .Z(r1164_n87) );
  EO r1164_U281 ( .A(r1164_n99), .B(r1164_n87), .Z(N2597) );
  IV r1164_U280 ( .A(U3_U6_Z_19), .Z(r1164_n82) );
  EO r1164_U279 ( .A(U3_U5_Z_19), .B(r1164_n82), .Z(r1164_n91) );
  NR2 r1164_U278 ( .A(U3_U5_Z_17), .B(r1164_n98), .Z(r1164_n96) );
  AO4 r1164_U277 ( .A(r1164_n94), .B(r1164_n95), .C(r1164_n96), .D(r1164_n97), 
        .Z(r1164_n92) );
  AN2 r1164_U276 ( .A(r1164_n92), .B(U3_U5_Z_18), .Z(r1164_n93) );
  AO4 r1164_U275 ( .A(U3_U5_Z_18), .B(r1164_n92), .C(U3_U6_Z_18), .D(r1164_n93), .Z(r1164_n80) );
  EO r1164_U274 ( .A(r1164_n91), .B(r1164_n80), .Z(N2598) );
  ND2 r1164_U273 ( .A(U3_U6_Z_0), .B(U3_U5_Z_0), .Z(r1164_n89) );
  EO r1164_U272 ( .A(U3_U6_Z_1), .B(U3_U5_Z_1), .Z(r1164_n90) );
  EN r1164_U271 ( .A(r1164_n89), .B(r1164_n90), .Z(N2580) );
  EN r1164_U270 ( .A(U3_U5_Z_20), .B(U3_U6_Z_20), .Z(r1164_n83) );
  IV r1164_U269 ( .A(U3_U5_Z_19), .Z(r1164_n79) );
  ND2 r1164_U268 ( .A(r1164_n87), .B(r1164_n88), .Z(r1164_n86) );
  EO1 r1164_U267 ( .A(r1164_n86), .B(U3_U6_Z_18), .C(r1164_n87), .D(r1164_n88), 
        .Z(r1164_n84) );
  OR2 r1164_U266 ( .A(r1164_n84), .B(r1164_n79), .Z(r1164_n85) );
  AO2 r1164_U265 ( .A(r1164_n79), .B(r1164_n84), .C(r1164_n82), .D(r1164_n85), 
        .Z(r1164_n74) );
  EN r1164_U264 ( .A(r1164_n83), .B(r1164_n74), .Z(N2599) );
  IV r1164_U263 ( .A(U3_U6_Z_21), .Z(r1164_n70) );
  EO r1164_U262 ( .A(U3_U5_Z_21), .B(r1164_n70), .Z(r1164_n76) );
  AN2 r1164_U261 ( .A(r1164_n80), .B(r1164_n79), .Z(r1164_n81) );
  AO4 r1164_U260 ( .A(r1164_n79), .B(r1164_n80), .C(r1164_n81), .D(r1164_n82), 
        .Z(r1164_n77) );
  AN2 r1164_U259 ( .A(r1164_n77), .B(U3_U5_Z_20), .Z(r1164_n78) );
  AO4 r1164_U258 ( .A(U3_U5_Z_20), .B(r1164_n77), .C(U3_U6_Z_20), .D(r1164_n78), .Z(r1164_n68) );
  EO r1164_U257 ( .A(r1164_n76), .B(r1164_n68), .Z(N2600) );
  EN r1164_U256 ( .A(U3_U5_Z_22), .B(U3_U6_Z_22), .Z(r1164_n71) );
  IV r1164_U255 ( .A(U3_U5_Z_21), .Z(r1164_n67) );
  OR2 r1164_U254 ( .A(r1164_n74), .B(U3_U5_Z_20), .Z(r1164_n75) );
  AO2 r1164_U253 ( .A(r1164_n74), .B(U3_U5_Z_20), .C(r1164_n75), .D(U3_U6_Z_20), .Z(r1164_n72) );
  OR2 r1164_U252 ( .A(r1164_n72), .B(r1164_n67), .Z(r1164_n73) );
  AO2 r1164_U251 ( .A(r1164_n67), .B(r1164_n72), .C(r1164_n70), .D(r1164_n73), 
        .Z(r1164_n62) );
  EN r1164_U250 ( .A(r1164_n71), .B(r1164_n62), .Z(N2601) );
  IV r1164_U249 ( .A(U3_U6_Z_23), .Z(r1164_n58) );
  EO r1164_U248 ( .A(U3_U5_Z_23), .B(r1164_n58), .Z(r1164_n64) );
  AN2 r1164_U247 ( .A(r1164_n68), .B(r1164_n67), .Z(r1164_n69) );
  AO4 r1164_U246 ( .A(r1164_n67), .B(r1164_n68), .C(r1164_n69), .D(r1164_n70), 
        .Z(r1164_n65) );
  AN2 r1164_U245 ( .A(r1164_n65), .B(U3_U5_Z_22), .Z(r1164_n66) );
  AO4 r1164_U244 ( .A(U3_U5_Z_22), .B(r1164_n65), .C(U3_U6_Z_22), .D(r1164_n66), .Z(r1164_n56) );
  EO r1164_U243 ( .A(r1164_n64), .B(r1164_n56), .Z(N2602) );
  EN r1164_U242 ( .A(U3_U5_Z_24), .B(U3_U6_Z_24), .Z(r1164_n59) );
  IV r1164_U241 ( .A(U3_U5_Z_23), .Z(r1164_n55) );
  OR2 r1164_U240 ( .A(r1164_n62), .B(U3_U5_Z_22), .Z(r1164_n63) );
  AO2 r1164_U239 ( .A(r1164_n62), .B(U3_U5_Z_22), .C(r1164_n63), .D(U3_U6_Z_22), .Z(r1164_n60) );
  OR2 r1164_U238 ( .A(r1164_n60), .B(r1164_n55), .Z(r1164_n61) );
  AO2 r1164_U237 ( .A(r1164_n55), .B(r1164_n60), .C(r1164_n58), .D(r1164_n61), 
        .Z(r1164_n51) );
  EN r1164_U236 ( .A(r1164_n59), .B(r1164_n51), .Z(N2603) );
  IV r1164_U235 ( .A(U3_U6_Z_25), .Z(r1164_n48) );
  EO r1164_U234 ( .A(U3_U5_Z_25), .B(r1164_n48), .Z(r1164_n52) );
  AN2 r1164_U233 ( .A(r1164_n56), .B(r1164_n55), .Z(r1164_n57) );
  AO4 r1164_U232 ( .A(r1164_n55), .B(r1164_n56), .C(r1164_n57), .D(r1164_n58), 
        .Z(r1164_n53) );
  AN2 r1164_U231 ( .A(r1164_n53), .B(U3_U5_Z_24), .Z(r1164_n54) );
  AO4 r1164_U230 ( .A(U3_U5_Z_24), .B(r1164_n53), .C(U3_U6_Z_24), .D(r1164_n54), .Z(r1164_n44) );
  EO r1164_U229 ( .A(r1164_n52), .B(r1164_n44), .Z(N2604) );
  IV r1164_U228 ( .A(U3_U6_Z_26), .Z(r1164_n38) );
  EO r1164_U227 ( .A(U3_U5_Z_26), .B(r1164_n38), .Z(r1164_n46) );
  IV r1164_U226 ( .A(U3_U5_Z_25), .Z(r1164_n43) );
  OR2 r1164_U225 ( .A(r1164_n51), .B(U3_U5_Z_24), .Z(r1164_n50) );
  AO2 r1164_U224 ( .A(r1164_n50), .B(U3_U6_Z_24), .C(r1164_n51), .D(U3_U5_Z_24), .Z(r1164_n47) );
  OR2 r1164_U223 ( .A(r1164_n47), .B(r1164_n43), .Z(r1164_n49) );
  AO2 r1164_U222 ( .A(r1164_n43), .B(r1164_n47), .C(r1164_n48), .D(r1164_n49), 
        .Z(r1164_n39) );
  EN r1164_U221 ( .A(r1164_n46), .B(r1164_n39), .Z(N2605) );
  EN r1164_U220 ( .A(U3_U5_Z_27), .B(U3_U6_Z_27), .Z(r1164_n40) );
  ND2 r1164_U219 ( .A(r1164_n44), .B(r1164_n43), .Z(r1164_n45) );
  EON1 r1164_U218 ( .A(r1164_n43), .B(r1164_n44), .C(r1164_n45), .D(U3_U6_Z_25), .Z(r1164_n42) );
  ND2 r1164_U217 ( .A(r1164_n42), .B(U3_U5_Z_26), .Z(r1164_n41) );
  EO1 r1164_U216 ( .A(r1164_n38), .B(r1164_n41), .C(U3_U5_Z_26), .D(r1164_n42), 
        .Z(r1164_n32) );
  EN r1164_U215 ( .A(r1164_n40), .B(r1164_n32), .Z(N2606) );
  IV r1164_U214 ( .A(U3_U6_Z_28), .Z(r1164_n25) );
  EO r1164_U213 ( .A(U3_U5_Z_28), .B(r1164_n25), .Z(r1164_n34) );
  NR2 r1164_U212 ( .A(r1164_n39), .B(U3_U5_Z_26), .Z(r1164_n37) );
  EON1 r1164_U211 ( .A(r1164_n37), .B(r1164_n38), .C(r1164_n39), .D(U3_U5_Z_26), .Z(r1164_n35) );
  AN2 r1164_U210 ( .A(r1164_n35), .B(U3_U5_Z_27), .Z(r1164_n36) );
  AO4 r1164_U209 ( .A(U3_U5_Z_27), .B(r1164_n35), .C(U3_U6_Z_27), .D(r1164_n36), .Z(r1164_n22) );
  EO r1164_U208 ( .A(r1164_n34), .B(r1164_n22), .Z(N2607) );
  EN r1164_U207 ( .A(U3_U6_Z_29), .B(U3_U5_Z_29), .Z(r1164_n28) );
  OR2 r1164_U206 ( .A(r1164_n32), .B(U3_U5_Z_27), .Z(r1164_n33) );
  AO2 r1164_U205 ( .A(U3_U5_Z_27), .B(r1164_n32), .C(r1164_n33), .D(U3_U6_Z_27), .Z(r1164_n31) );
  IV r1164_U204 ( .A(U3_U5_Z_28), .Z(r1164_n23) );
  NR2 r1164_U203 ( .A(r1164_n31), .B(r1164_n23), .Z(r1164_n30) );
  EON1 r1164_U202 ( .A(U3_U6_Z_28), .B(r1164_n30), .C(r1164_n23), .D(r1164_n31), .Z(r1164_n29) );
  EO r1164_U201 ( .A(r1164_n28), .B(r1164_n29), .Z(N2608) );
  EN r1164_U200 ( .A(U3_U6_Z_2), .B(U3_U5_Z_2), .Z(r1164_n26) );
  EO r1164_U199 ( .A(r1164_n26), .B(r1164_n27), .Z(N2581) );
  EN r1164_U198 ( .A(U3_U6_Z_30), .B(U3_U5_Z_30), .Z(r1164_n18) );
  AN2 r1164_U197 ( .A(r1164_n22), .B(r1164_n23), .Z(r1164_n24) );
  AO4 r1164_U196 ( .A(r1164_n22), .B(r1164_n23), .C(r1164_n24), .D(r1164_n25), 
        .Z(r1164_n20) );
  AN2 r1164_U195 ( .A(r1164_n20), .B(U3_U5_Z_29), .Z(r1164_n21) );
  AO4 r1164_U194 ( .A(U3_U5_Z_29), .B(r1164_n20), .C(U3_U6_Z_29), .D(r1164_n21), .Z(r1164_n19) );
  EO r1164_U193 ( .A(r1164_n18), .B(r1164_n19), .Z(N2609) );
  EN r1164_U192 ( .A(U3_U6_Z_3), .B(U3_U5_Z_3), .Z(r1164_n17) );
  EO r1164_U191 ( .A(r1164_n16), .B(r1164_n17), .Z(N2582) );
  EN r1164_U190 ( .A(U3_U6_Z_4), .B(U3_U5_Z_4), .Z(r1164_n15) );
  EO r1164_U189 ( .A(r1164_n14), .B(r1164_n15), .Z(N2583) );
  EN r1164_U188 ( .A(U3_U6_Z_5), .B(U3_U5_Z_5), .Z(r1164_n12) );
  EO r1164_U187 ( .A(r1164_n12), .B(r1164_n13), .Z(N2584) );
  EN r1164_U186 ( .A(U3_U6_Z_6), .B(U3_U5_Z_6), .Z(r1164_n11) );
  EO r1164_U185 ( .A(r1164_n10), .B(r1164_n11), .Z(N2585) );
  EN r1164_U184 ( .A(U3_U6_Z_7), .B(U3_U5_Z_7), .Z(r1164_n8) );
  EO r1164_U183 ( .A(r1164_n8), .B(r1164_n9), .Z(N2586) );
  EO r1164_U182 ( .A(U3_U6_Z_8), .B(r1164_n6), .Z(r1164_n7) );
  EO r1164_U181 ( .A(r1164_n5), .B(r1164_n7), .Z(N2587) );
  EN r1164_U180 ( .A(U3_U6_Z_9), .B(U3_U5_Z_9), .Z(r1164_n1) );
  NR2 r1164_U179 ( .A(r1164_n5), .B(r1164_n6), .Z(r1164_n4) );
  AO4 r1164_U178 ( .A(U3_U5_Z_8), .B(r1164_n3), .C(U3_U6_Z_8), .D(r1164_n4), 
        .Z(r1164_n2) );
  EO r1164_U177 ( .A(r1164_n1), .B(r1164_n2), .Z(N2588) );
  EO r1166_U274 ( .A(U3_U22_Z_0), .B(U3_U23_Z_0), .Z(r1166_n106) );
  EO r1166_U273 ( .A(U3_U21_Z_0), .B(U3_U23_Z_0), .Z(r1166_n107) );
  EO r1166_U272 ( .A(r1166_n106), .B(r1166_n107), .Z(n234) );
  IV r1166_U271 ( .A(U3_U23_Z_0), .Z(r1166_n27) );
  EN r1166_U270 ( .A(U3_U22_Z_10), .B(r1166_n27), .Z(r1166_n103) );
  EO r1166_U269 ( .A(U3_U22_Z_7), .B(U3_U23_Z_0), .Z(r1166_n6) );
  EN r1166_U268 ( .A(U3_U22_Z_8), .B(r1166_n27), .Z(r1166_n3) );
  EO r1166_U267 ( .A(U3_U22_Z_5), .B(U3_U23_Z_0), .Z(r1166_n10) );
  EN r1166_U266 ( .A(U3_U22_Z_6), .B(r1166_n27), .Z(r1166_n7) );
  EO r1166_U265 ( .A(U3_U22_Z_3), .B(r1166_n27), .Z(r1166_n15) );
  IV r1166_U264 ( .A(r1166_n15), .Z(r1166_n14) );
  EO r1166_U263 ( .A(U3_U22_Z_4), .B(r1166_n27), .Z(r1166_n11) );
  IV r1166_U262 ( .A(r1166_n11), .Z(r1166_n105) );
  EN r1166_U261 ( .A(U3_U22_Z_2), .B(U3_U23_Z_0), .Z(r1166_n32) );
  EO r1166_U260 ( .A(U3_U22_Z_1), .B(r1166_n27), .Z(r1166_n33) );
  AO5 r1166_U259 ( .A(U3_U23_Z_0), .B(U3_U21_Z_0), .C(r1166_n106), .Z(
        r1166_n34) );
  OR3 r1166_U258 ( .A(r1166_n32), .B(r1166_n33), .C(r1166_n34), .Z(r1166_n16)
         );
  IV r1166_U257 ( .A(r1166_n16), .Z(r1166_n13) );
  AN3 r1166_U256 ( .A(r1166_n14), .B(r1166_n105), .C(r1166_n13), .Z(r1166_n9)
         );
  AN3 r1166_U255 ( .A(r1166_n10), .B(r1166_n7), .C(r1166_n9), .Z(r1166_n5) );
  AN3 r1166_U254 ( .A(r1166_n6), .B(r1166_n3), .C(r1166_n5), .Z(r1166_n2) );
  EN r1166_U253 ( .A(U3_U22_Z_9), .B(r1166_n27), .Z(r1166_n1) );
  ND2 r1166_U252 ( .A(r1166_n2), .B(r1166_n1), .Z(r1166_n104) );
  EN r1166_U251 ( .A(r1166_n103), .B(r1166_n104), .Z(n224) );
  EO r1166_U250 ( .A(U3_U22_Z_11), .B(r1166_n27), .Z(r1166_n101) );
  ND3 r1166_U249 ( .A(r1166_n103), .B(r1166_n1), .C(r1166_n2), .Z(r1166_n102)
         );
  EO r1166_U248 ( .A(r1166_n101), .B(r1166_n102), .Z(n223) );
  EO r1166_U247 ( .A(U3_U22_Z_12), .B(r1166_n27), .Z(r1166_n99) );
  IV r1166_U246 ( .A(r1166_n102), .Z(r1166_n98) );
  IV r1166_U245 ( .A(r1166_n101), .Z(r1166_n97) );
  ND2 r1166_U244 ( .A(r1166_n98), .B(r1166_n97), .Z(r1166_n100) );
  EO r1166_U243 ( .A(r1166_n99), .B(r1166_n100), .Z(n222) );
  EO r1166_U242 ( .A(U3_U22_Z_13), .B(U3_U23_Z_0), .Z(r1166_n92) );
  IV r1166_U241 ( .A(r1166_n99), .Z(r1166_n96) );
  AN3 r1166_U240 ( .A(r1166_n96), .B(r1166_n97), .C(r1166_n98), .Z(r1166_n94)
         );
  EO r1166_U239 ( .A(r1166_n92), .B(r1166_n94), .Z(n221) );
  EN r1166_U238 ( .A(U3_U22_Z_14), .B(r1166_n27), .Z(r1166_n93) );
  ND2 r1166_U237 ( .A(r1166_n94), .B(r1166_n92), .Z(r1166_n95) );
  EN r1166_U236 ( .A(r1166_n93), .B(r1166_n95), .Z(n220) );
  EO r1166_U235 ( .A(U3_U22_Z_15), .B(r1166_n27), .Z(r1166_n90) );
  ND3 r1166_U234 ( .A(r1166_n92), .B(r1166_n93), .C(r1166_n94), .Z(r1166_n91)
         );
  EO r1166_U233 ( .A(r1166_n90), .B(r1166_n91), .Z(n219) );
  EN r1166_U232 ( .A(n2141), .B(r1166_n27), .Z(r1166_n84) );
  NR2 r1166_U231 ( .A(r1166_n90), .B(r1166_n91), .Z(r1166_n85) );
  EO r1166_U230 ( .A(r1166_n85), .B(U3_U21_Z_16), .Z(r1166_n89) );
  EO r1166_U229 ( .A(r1166_n84), .B(r1166_n89), .Z(n218) );
  EO r1166_U228 ( .A(n2142), .B(U3_U23_Z_0), .Z(r1166_n81) );
  EO r1166_U227 ( .A(n2141), .B(U3_U23_Z_0), .Z(r1166_n88) );
  AO5 r1166_U226 ( .A(r1166_n85), .B(U3_U21_Z_16), .C(r1166_n88), .Z(r1166_n87) );
  EN r1166_U225 ( .A(r1166_n87), .B(U3_U21_Z_17), .Z(r1166_n86) );
  EO r1166_U224 ( .A(r1166_n81), .B(r1166_n86), .Z(n217) );
  EO r1166_U223 ( .A(n2143), .B(r1166_n27), .Z(r1166_n77) );
  ND2 r1166_U222 ( .A(r1166_n85), .B(r1166_n84), .Z(r1166_n82) );
  IV r1166_U221 ( .A(U3_U21_Z_16), .Z(r1166_n83) );
  EO1 r1166_U220 ( .A(r1166_n82), .B(r1166_n83), .C(r1166_n84), .D(r1166_n85), 
        .Z(r1166_n80) );
  AO5 r1166_U219 ( .A(r1166_n80), .B(U3_U21_Z_17), .C(r1166_n81), .Z(r1166_n78) );
  EN r1166_U218 ( .A(r1166_n78), .B(U3_U21_Z_18), .Z(r1166_n79) );
  EN r1166_U217 ( .A(r1166_n77), .B(r1166_n79), .Z(n216) );
  EO r1166_U216 ( .A(n2144), .B(r1166_n27), .Z(r1166_n72) );
  ND2 r1166_U215 ( .A(r1166_n78), .B(r1166_n77), .Z(r1166_n76) );
  EO1 r1166_U214 ( .A(r1166_n76), .B(U3_U21_Z_18), .C(r1166_n77), .D(r1166_n78), .Z(r1166_n73) );
  EN r1166_U213 ( .A(r1166_n73), .B(U3_U21_Z_19), .Z(r1166_n75) );
  EN r1166_U212 ( .A(r1166_n72), .B(r1166_n75), .Z(n215) );
  EO r1166_U211 ( .A(r1166_n33), .B(r1166_n34), .Z(n233) );
  EN r1166_U210 ( .A(U3_U22_Z_20), .B(r1166_n27), .Z(r1166_n68) );
  NR2 r1166_U209 ( .A(r1166_n73), .B(r1166_n72), .Z(r1166_n74) );
  EO1 r1166_U208 ( .A(r1166_n72), .B(r1166_n73), .C(U3_U21_Z_19), .D(r1166_n74), .Z(r1166_n69) );
  EO r1166_U207 ( .A(r1166_n69), .B(U3_U21_Z_20), .Z(r1166_n71) );
  EO r1166_U206 ( .A(r1166_n68), .B(r1166_n71), .Z(n214) );
  EO r1166_U205 ( .A(U3_U22_Z_21), .B(r1166_n27), .Z(r1166_n64) );
  OR2 r1166_U204 ( .A(r1166_n69), .B(r1166_n68), .Z(r1166_n70) );
  AO2 r1166_U203 ( .A(r1166_n68), .B(r1166_n69), .C(r1166_n70), .D(U3_U21_Z_20), .Z(r1166_n65) );
  EN r1166_U202 ( .A(r1166_n65), .B(U3_U21_Z_21), .Z(r1166_n67) );
  EN r1166_U201 ( .A(r1166_n64), .B(r1166_n67), .Z(n213) );
  EN r1166_U200 ( .A(U3_U22_Z_22), .B(r1166_n27), .Z(r1166_n60) );
  NR2 r1166_U199 ( .A(r1166_n65), .B(r1166_n64), .Z(r1166_n66) );
  EO1 r1166_U198 ( .A(r1166_n64), .B(r1166_n65), .C(U3_U21_Z_21), .D(r1166_n66), .Z(r1166_n61) );
  EO r1166_U197 ( .A(r1166_n61), .B(U3_U21_Z_22), .Z(r1166_n63) );
  EO r1166_U196 ( .A(r1166_n60), .B(r1166_n63), .Z(n212) );
  EO r1166_U195 ( .A(U3_U22_Z_23), .B(r1166_n27), .Z(r1166_n56) );
  OR2 r1166_U194 ( .A(r1166_n61), .B(r1166_n60), .Z(r1166_n62) );
  AO2 r1166_U193 ( .A(r1166_n60), .B(r1166_n61), .C(r1166_n62), .D(U3_U21_Z_22), .Z(r1166_n57) );
  EN r1166_U192 ( .A(r1166_n57), .B(U3_U21_Z_23), .Z(r1166_n59) );
  EN r1166_U191 ( .A(r1166_n56), .B(r1166_n59), .Z(n211) );
  EN r1166_U190 ( .A(U3_U22_Z_24), .B(r1166_n27), .Z(r1166_n52) );
  NR2 r1166_U189 ( .A(r1166_n57), .B(r1166_n56), .Z(r1166_n58) );
  EO1 r1166_U188 ( .A(r1166_n56), .B(r1166_n57), .C(U3_U21_Z_23), .D(r1166_n58), .Z(r1166_n53) );
  EO r1166_U187 ( .A(r1166_n53), .B(U3_U21_Z_24), .Z(r1166_n55) );
  EO r1166_U186 ( .A(r1166_n52), .B(r1166_n55), .Z(n210) );
  EO r1166_U185 ( .A(U3_U22_Z_25), .B(r1166_n27), .Z(r1166_n48) );
  OR2 r1166_U184 ( .A(r1166_n53), .B(r1166_n52), .Z(r1166_n54) );
  AO2 r1166_U183 ( .A(r1166_n52), .B(r1166_n53), .C(r1166_n54), .D(U3_U21_Z_24), .Z(r1166_n49) );
  EN r1166_U182 ( .A(r1166_n49), .B(U3_U21_Z_25), .Z(r1166_n51) );
  EN r1166_U181 ( .A(r1166_n48), .B(r1166_n51), .Z(n209) );
  EN r1166_U180 ( .A(U3_U22_Z_26), .B(r1166_n27), .Z(r1166_n44) );
  NR2 r1166_U179 ( .A(r1166_n49), .B(r1166_n48), .Z(r1166_n50) );
  EO1 r1166_U178 ( .A(r1166_n48), .B(r1166_n49), .C(U3_U21_Z_25), .D(r1166_n50), .Z(r1166_n45) );
  EO r1166_U177 ( .A(r1166_n45), .B(U3_U21_Z_26), .Z(r1166_n47) );
  EO r1166_U176 ( .A(r1166_n44), .B(r1166_n47), .Z(n208) );
  EO r1166_U175 ( .A(U3_U22_Z_27), .B(r1166_n27), .Z(r1166_n40) );
  OR2 r1166_U174 ( .A(r1166_n45), .B(r1166_n44), .Z(r1166_n46) );
  AO2 r1166_U173 ( .A(r1166_n44), .B(r1166_n45), .C(r1166_n46), .D(U3_U21_Z_26), .Z(r1166_n41) );
  EN r1166_U172 ( .A(r1166_n41), .B(U3_U21_Z_27), .Z(r1166_n43) );
  EN r1166_U171 ( .A(r1166_n40), .B(r1166_n43), .Z(n207) );
  EN r1166_U170 ( .A(U3_U22_Z_28), .B(r1166_n27), .Z(r1166_n36) );
  NR2 r1166_U169 ( .A(r1166_n41), .B(r1166_n40), .Z(r1166_n42) );
  EO1 r1166_U168 ( .A(r1166_n40), .B(r1166_n41), .C(U3_U21_Z_27), .D(r1166_n42), .Z(r1166_n37) );
  EO r1166_U167 ( .A(r1166_n37), .B(U3_U21_Z_28), .Z(r1166_n39) );
  EO r1166_U166 ( .A(r1166_n36), .B(r1166_n39), .Z(n206) );
  EO r1166_U165 ( .A(U3_U22_Z_29), .B(r1166_n27), .Z(r1166_n24) );
  IV r1166_U164 ( .A(r1166_n24), .Z(r1166_n25) );
  OR2 r1166_U163 ( .A(r1166_n37), .B(r1166_n36), .Z(r1166_n38) );
  AO2 r1166_U162 ( .A(r1166_n36), .B(r1166_n37), .C(r1166_n38), .D(U3_U21_Z_28), .Z(r1166_n23) );
  IV r1166_U161 ( .A(U3_U21_Z_29), .Z(r1166_n22) );
  EO r1166_U160 ( .A(r1166_n23), .B(r1166_n22), .Z(r1166_n35) );
  EO r1166_U159 ( .A(r1166_n25), .B(r1166_n35), .Z(n205) );
  NR2 r1166_U158 ( .A(r1166_n33), .B(r1166_n34), .Z(r1166_n31) );
  EN r1166_U157 ( .A(r1166_n31), .B(r1166_n32), .Z(n232) );
  EO r1166_U156 ( .A(U3_U22_Z_30), .B(U3_U23_Z_0), .Z(r1166_n20) );
  IV r1166_U155 ( .A(r1166_n23), .Z(r1166_n26) );
  NR2 r1166_U154 ( .A(r1166_n23), .B(r1166_n24), .Z(r1166_n30) );
  AO4 r1166_U153 ( .A(r1166_n25), .B(r1166_n26), .C(U3_U21_Z_29), .D(r1166_n30), .Z(r1166_n29) );
  EN r1166_U152 ( .A(r1166_n29), .B(U3_U21_Z_30), .Z(r1166_n28) );
  EO r1166_U151 ( .A(r1166_n20), .B(r1166_n28), .Z(n204) );
  EO r1166_U150 ( .A(U3_U22_Z_31), .B(r1166_n27), .Z(r1166_n17) );
  ND2 r1166_U149 ( .A(r1166_n25), .B(r1166_n26), .Z(r1166_n21) );
  AO2 r1166_U148 ( .A(r1166_n21), .B(r1166_n22), .C(r1166_n23), .D(r1166_n24), 
        .Z(r1166_n19) );
  AO5 r1166_U147 ( .A(r1166_n19), .B(U3_U21_Z_30), .C(r1166_n20), .Z(r1166_n18) );
  EO r1166_U146 ( .A(r1166_n17), .B(r1166_n18), .Z(n203) );
  EO r1166_U145 ( .A(r1166_n15), .B(r1166_n16), .Z(n231) );
  ND2 r1166_U144 ( .A(r1166_n13), .B(r1166_n14), .Z(r1166_n12) );
  EO r1166_U143 ( .A(r1166_n11), .B(r1166_n12), .Z(n230) );
  EO r1166_U142 ( .A(r1166_n10), .B(r1166_n9), .Z(n229) );
  ND2 r1166_U141 ( .A(r1166_n9), .B(r1166_n10), .Z(r1166_n8) );
  EN r1166_U140 ( .A(r1166_n7), .B(r1166_n8), .Z(n228) );
  EO r1166_U139 ( .A(r1166_n6), .B(r1166_n5), .Z(n227) );
  ND2 r1166_U138 ( .A(r1166_n5), .B(r1166_n6), .Z(r1166_n4) );
  EN r1166_U137 ( .A(r1166_n3), .B(r1166_n4), .Z(n226) );
  EO r1166_U136 ( .A(r1166_n1), .B(r1166_n2), .Z(n225) );
  EO r253_U344 ( .A(U3_U14_Z_7), .B(U3_U19_Z_0), .Z(r253_n49) );
  EO r253_U343 ( .A(U3_U18_Z_0), .B(U3_U14_Z_7), .Z(r253_n148) );
  EO r253_U342 ( .A(r253_n49), .B(r253_n148), .Z(n317) );
  IV r253_U341 ( .A(U3_U14_Z_7), .Z(r253_n37) );
  EO r253_U340 ( .A(r253_n37), .B(U3_U18_Z_10), .Z(r253_n135) );
  EO r253_U339 ( .A(U3_U19_Z_7), .B(r253_n37), .Z(r253_n7) );
  EN r253_U338 ( .A(U3_U19_Z_6), .B(r253_n37), .Z(r253_n10) );
  EO r253_U337 ( .A(U3_U19_Z_5), .B(r253_n37), .Z(r253_n23) );
  EN r253_U336 ( .A(U3_U19_Z_3), .B(r253_n37), .Z(r253_n25) );
  IV r253_U335 ( .A(U3_U18_Z_2), .Z(r253_n31) );
  EN r253_U334 ( .A(n5490), .B(r253_n37), .Z(r253_n94) );
  NR2 r253_U333 ( .A(r253_n94), .B(U3_U18_Z_1), .Z(r253_n48) );
  MUX21L r253_U332 ( .A(U3_U14_Z_7), .B(U3_U18_Z_0), .S(U3_U19_Z_0), .Z(
        r253_n93) );
  ND2 r253_U331 ( .A(U3_U18_Z_1), .B(r253_n94), .Z(r253_n95) );
  AO7 r253_U330 ( .A(r253_n48), .B(r253_n93), .C(r253_n95), .Z(r253_n147) );
  EO r253_U329 ( .A(U3_U19_Z_2), .B(r253_n37), .Z(r253_n29) );
  IV r253_U328 ( .A(r253_n29), .Z(r253_n42) );
  ND2 r253_U327 ( .A(r253_n147), .B(r253_n42), .Z(r253_n146) );
  EO1 r253_U326 ( .A(r253_n31), .B(r253_n146), .C(r253_n42), .D(r253_n147), 
        .Z(r253_n33) );
  OR2 r253_U325 ( .A(r253_n33), .B(r253_n25), .Z(r253_n145) );
  AO2 r253_U324 ( .A(r253_n25), .B(r253_n33), .C(r253_n145), .D(U3_U18_Z_3), 
        .Z(r253_n144) );
  EO r253_U323 ( .A(U3_U19_Z_4), .B(r253_n37), .Z(r253_n16) );
  NR2 r253_U322 ( .A(r253_n144), .B(r253_n16), .Z(r253_n143) );
  EON1 r253_U321 ( .A(U3_U18_Z_4), .B(r253_n143), .C(r253_n16), .D(r253_n144), 
        .Z(r253_n21) );
  AN2 r253_U320 ( .A(r253_n21), .B(r253_n23), .Z(r253_n142) );
  IV r253_U319 ( .A(U3_U18_Z_5), .Z(r253_n22) );
  AO4 r253_U318 ( .A(r253_n23), .B(r253_n21), .C(r253_n142), .D(r253_n22), .Z(
        r253_n140) );
  AN2 r253_U317 ( .A(r253_n140), .B(r253_n10), .Z(r253_n141) );
  AO4 r253_U316 ( .A(r253_n10), .B(r253_n140), .C(U3_U18_Z_6), .D(r253_n141), 
        .Z(r253_n9) );
  ND2 r253_U315 ( .A(r253_n9), .B(r253_n7), .Z(r253_n139) );
  EON1 r253_U314 ( .A(r253_n7), .B(r253_n9), .C(r253_n139), .D(U3_U18_Z_7), 
        .Z(r253_n133) );
  ND2 r253_U313 ( .A(U3_U14_Z_7), .B(r253_n133), .Z(r253_n138) );
  IV r253_U312 ( .A(U3_U18_Z_8), .Z(r253_n6) );
  IV r253_U311 ( .A(r253_n133), .Z(r253_n4) );
  AO2 r253_U310 ( .A(r253_n138), .B(r253_n6), .C(r253_n4), .D(r253_n37), .Z(
        r253_n137) );
  AO5 r253_U309 ( .A(U3_U14_Z_7), .B(U3_U18_Z_9), .C(r253_n137), .Z(r253_n136)
         );
  EO r253_U308 ( .A(r253_n135), .B(r253_n136), .Z(n307) );
  EO r253_U307 ( .A(r253_n37), .B(U3_U18_Z_11), .Z(r253_n130) );
  NR2 r253_U306 ( .A(r253_n4), .B(r253_n37), .Z(r253_n134) );
  AO4 r253_U305 ( .A(U3_U14_Z_7), .B(r253_n133), .C(U3_U18_Z_8), .D(r253_n134), 
        .Z(r253_n2) );
  OR2 r253_U304 ( .A(r253_n2), .B(r253_n37), .Z(r253_n132) );
  IV r253_U303 ( .A(U3_U18_Z_9), .Z(r253_n3) );
  AO2 r253_U302 ( .A(r253_n132), .B(r253_n3), .C(r253_n2), .D(r253_n37), .Z(
        r253_n131) );
  AO5 r253_U301 ( .A(U3_U14_Z_7), .B(U3_U18_Z_10), .C(r253_n131), .Z(r253_n129) );
  EO r253_U300 ( .A(r253_n130), .B(r253_n129), .Z(n306) );
  ND2 r253_U299 ( .A(r253_n129), .B(r253_n37), .Z(r253_n128) );
  EO1 r253_U298 ( .A(r253_n128), .B(U3_U18_Z_11), .C(r253_n37), .D(r253_n129), 
        .Z(r253_n123) );
  IV r253_U297 ( .A(U3_U18_Z_12), .Z(r253_n122) );
  EO r253_U296 ( .A(U3_U14_Z_7), .B(r253_n122), .Z(r253_n127) );
  EO r253_U295 ( .A(r253_n123), .B(r253_n127), .Z(n305) );
  IV r253_U294 ( .A(U3_U18_Z_13), .Z(r253_n116) );
  EO r253_U293 ( .A(U3_U14_Z_7), .B(r253_n116), .Z(r253_n125) );
  IV r253_U292 ( .A(r253_n123), .Z(r253_n124) );
  NR2 r253_U291 ( .A(r253_n123), .B(r253_n37), .Z(r253_n126) );
  AO4 r253_U290 ( .A(U3_U14_Z_7), .B(r253_n124), .C(U3_U18_Z_12), .D(r253_n126), .Z(r253_n117) );
  EO r253_U289 ( .A(r253_n125), .B(r253_n117), .Z(n304) );
  EO r253_U288 ( .A(r253_n37), .B(U3_U18_Z_14), .Z(r253_n118) );
  ND2 r253_U287 ( .A(U3_U14_Z_7), .B(r253_n124), .Z(r253_n121) );
  AO2 r253_U286 ( .A(r253_n121), .B(r253_n122), .C(r253_n123), .D(r253_n37), 
        .Z(r253_n120) );
  AO5 r253_U285 ( .A(U3_U14_Z_7), .B(U3_U18_Z_13), .C(r253_n120), .Z(r253_n119) );
  EO r253_U284 ( .A(r253_n118), .B(r253_n119), .Z(n303) );
  EO r253_U283 ( .A(r253_n37), .B(U3_U18_Z_15), .Z(r253_n113) );
  OR2 r253_U282 ( .A(r253_n117), .B(r253_n37), .Z(r253_n115) );
  AO2 r253_U281 ( .A(r253_n115), .B(r253_n116), .C(r253_n117), .D(r253_n37), 
        .Z(r253_n114) );
  AO5 r253_U280 ( .A(U3_U14_Z_7), .B(U3_U18_Z_14), .C(r253_n114), .Z(r253_n112) );
  EO r253_U279 ( .A(r253_n113), .B(r253_n112), .Z(n302) );
  ND2 r253_U278 ( .A(r253_n112), .B(r253_n37), .Z(r253_n111) );
  EO1 r253_U277 ( .A(r253_n111), .B(U3_U18_Z_15), .C(r253_n37), .D(r253_n112), 
        .Z(r253_n106) );
  IV r253_U276 ( .A(U3_U18_Z_16), .Z(r253_n105) );
  EO r253_U275 ( .A(U3_U14_Z_7), .B(r253_n105), .Z(r253_n110) );
  EO r253_U274 ( .A(r253_n106), .B(r253_n110), .Z(n301) );
  IV r253_U273 ( .A(U3_U18_Z_17), .Z(r253_n99) );
  EO r253_U272 ( .A(U3_U14_Z_7), .B(r253_n99), .Z(r253_n108) );
  IV r253_U271 ( .A(r253_n106), .Z(r253_n107) );
  NR2 r253_U270 ( .A(r253_n106), .B(r253_n37), .Z(r253_n109) );
  AO4 r253_U269 ( .A(U3_U14_Z_7), .B(r253_n107), .C(U3_U18_Z_16), .D(r253_n109), .Z(r253_n100) );
  EO r253_U268 ( .A(r253_n108), .B(r253_n100), .Z(n300) );
  EO r253_U267 ( .A(r253_n37), .B(U3_U18_Z_18), .Z(r253_n101) );
  ND2 r253_U266 ( .A(U3_U14_Z_7), .B(r253_n107), .Z(r253_n104) );
  AO2 r253_U265 ( .A(r253_n104), .B(r253_n105), .C(r253_n106), .D(r253_n37), 
        .Z(r253_n103) );
  AO5 r253_U264 ( .A(U3_U14_Z_7), .B(U3_U18_Z_17), .C(r253_n103), .Z(r253_n102) );
  EO r253_U263 ( .A(r253_n101), .B(r253_n102), .Z(n299) );
  EO r253_U262 ( .A(r253_n37), .B(U3_U18_Z_19), .Z(r253_n96) );
  OR2 r253_U261 ( .A(r253_n100), .B(r253_n37), .Z(r253_n98) );
  AO2 r253_U260 ( .A(r253_n98), .B(r253_n99), .C(r253_n100), .D(r253_n37), .Z(
        r253_n97) );
  AO5 r253_U259 ( .A(U3_U14_Z_7), .B(U3_U18_Z_18), .C(r253_n97), .Z(r253_n90)
         );
  EO r253_U258 ( .A(r253_n96), .B(r253_n90), .Z(n298) );
  IV r253_U257 ( .A(r253_n95), .Z(r253_n44) );
  NR2 r253_U256 ( .A(r253_n44), .B(r253_n48), .Z(r253_n91) );
  EN r253_U255 ( .A(r253_n94), .B(U3_U18_Z_1), .Z(r253_n92) );
  MUX21L r253_U254 ( .A(r253_n91), .B(r253_n92), .S(r253_n93), .Z(n316) );
  ND2 r253_U253 ( .A(r253_n90), .B(r253_n37), .Z(r253_n89) );
  EO1 r253_U252 ( .A(r253_n89), .B(U3_U18_Z_19), .C(r253_n37), .D(r253_n90), 
        .Z(r253_n84) );
  IV r253_U251 ( .A(U3_U18_Z_20), .Z(r253_n83) );
  EO r253_U250 ( .A(U3_U14_Z_7), .B(r253_n83), .Z(r253_n88) );
  EO r253_U249 ( .A(r253_n84), .B(r253_n88), .Z(n297) );
  IV r253_U248 ( .A(U3_U18_Z_21), .Z(r253_n77) );
  EO r253_U247 ( .A(U3_U14_Z_7), .B(r253_n77), .Z(r253_n86) );
  IV r253_U246 ( .A(r253_n84), .Z(r253_n85) );
  NR2 r253_U245 ( .A(r253_n84), .B(r253_n37), .Z(r253_n87) );
  AO4 r253_U244 ( .A(U3_U14_Z_7), .B(r253_n85), .C(U3_U18_Z_20), .D(r253_n87), 
        .Z(r253_n78) );
  EO r253_U243 ( .A(r253_n86), .B(r253_n78), .Z(n296) );
  EO r253_U242 ( .A(r253_n37), .B(U3_U18_Z_22), .Z(r253_n79) );
  ND2 r253_U241 ( .A(U3_U14_Z_7), .B(r253_n85), .Z(r253_n82) );
  AO2 r253_U240 ( .A(r253_n82), .B(r253_n83), .C(r253_n84), .D(r253_n37), .Z(
        r253_n81) );
  AO5 r253_U239 ( .A(U3_U14_Z_7), .B(U3_U18_Z_21), .C(r253_n81), .Z(r253_n80)
         );
  EO r253_U238 ( .A(r253_n79), .B(r253_n80), .Z(n295) );
  EO r253_U237 ( .A(r253_n37), .B(U3_U18_Z_23), .Z(r253_n74) );
  OR2 r253_U236 ( .A(r253_n78), .B(r253_n37), .Z(r253_n76) );
  AO2 r253_U235 ( .A(r253_n76), .B(r253_n77), .C(r253_n78), .D(r253_n37), .Z(
        r253_n75) );
  AO5 r253_U234 ( .A(U3_U14_Z_7), .B(U3_U18_Z_22), .C(r253_n75), .Z(r253_n73)
         );
  EO r253_U233 ( .A(r253_n74), .B(r253_n73), .Z(n294) );
  ND2 r253_U232 ( .A(r253_n73), .B(r253_n37), .Z(r253_n72) );
  EO1 r253_U231 ( .A(r253_n72), .B(U3_U18_Z_23), .C(r253_n37), .D(r253_n73), 
        .Z(r253_n67) );
  IV r253_U230 ( .A(U3_U18_Z_24), .Z(r253_n66) );
  EO r253_U229 ( .A(U3_U14_Z_7), .B(r253_n66), .Z(r253_n71) );
  EO r253_U228 ( .A(r253_n67), .B(r253_n71), .Z(n293) );
  IV r253_U227 ( .A(U3_U18_Z_25), .Z(r253_n60) );
  EO r253_U226 ( .A(U3_U14_Z_7), .B(r253_n60), .Z(r253_n69) );
  IV r253_U225 ( .A(r253_n67), .Z(r253_n68) );
  NR2 r253_U224 ( .A(r253_n67), .B(r253_n37), .Z(r253_n70) );
  AO4 r253_U223 ( .A(U3_U14_Z_7), .B(r253_n68), .C(U3_U18_Z_24), .D(r253_n70), 
        .Z(r253_n61) );
  EO r253_U222 ( .A(r253_n69), .B(r253_n61), .Z(n292) );
  EO r253_U221 ( .A(r253_n37), .B(U3_U18_Z_26), .Z(r253_n62) );
  ND2 r253_U220 ( .A(U3_U14_Z_7), .B(r253_n68), .Z(r253_n65) );
  AO2 r253_U219 ( .A(r253_n65), .B(r253_n66), .C(r253_n67), .D(r253_n37), .Z(
        r253_n64) );
  AO5 r253_U218 ( .A(U3_U14_Z_7), .B(U3_U18_Z_25), .C(r253_n64), .Z(r253_n63)
         );
  EO r253_U217 ( .A(r253_n62), .B(r253_n63), .Z(n291) );
  EO r253_U216 ( .A(r253_n37), .B(U3_U18_Z_27), .Z(r253_n57) );
  OR2 r253_U215 ( .A(r253_n61), .B(r253_n37), .Z(r253_n59) );
  AO2 r253_U214 ( .A(r253_n59), .B(r253_n60), .C(r253_n61), .D(r253_n37), .Z(
        r253_n58) );
  AO5 r253_U213 ( .A(U3_U14_Z_7), .B(U3_U18_Z_26), .C(r253_n58), .Z(r253_n56)
         );
  EO r253_U212 ( .A(r253_n57), .B(r253_n56), .Z(n290) );
  ND2 r253_U211 ( .A(r253_n56), .B(r253_n37), .Z(r253_n55) );
  EO1 r253_U210 ( .A(r253_n55), .B(U3_U18_Z_27), .C(r253_n37), .D(r253_n56), 
        .Z(r253_n51) );
  IV r253_U209 ( .A(U3_U18_Z_28), .Z(r253_n52) );
  EO r253_U208 ( .A(U3_U14_Z_7), .B(r253_n52), .Z(r253_n54) );
  EO r253_U207 ( .A(r253_n51), .B(r253_n54), .Z(n289) );
  EO r253_U206 ( .A(r253_n37), .B(U3_U18_Z_29), .Z(r253_n50) );
  OR2 r253_U205 ( .A(r253_n51), .B(r253_n37), .Z(r253_n53) );
  AO2 r253_U204 ( .A(r253_n37), .B(r253_n51), .C(r253_n52), .D(r253_n53), .Z(
        r253_n40) );
  EN r253_U203 ( .A(r253_n50), .B(r253_n40), .Z(n288) );
  IV r253_U202 ( .A(r253_n49), .Z(r253_n46) );
  AO6 r253_U201 ( .A(r253_n49), .B(U3_U14_Z_7), .C(U3_U18_Z_0), .Z(r253_n47)
         );
  AO1 r253_U200 ( .A(r253_n37), .B(r253_n46), .C(r253_n47), .D(r253_n48), .Z(
        r253_n45) );
  NR2 r253_U199 ( .A(r253_n44), .B(r253_n45), .Z(r253_n28) );
  EO r253_U198 ( .A(r253_n28), .B(r253_n31), .Z(r253_n43) );
  EO r253_U197 ( .A(r253_n42), .B(r253_n43), .Z(n315) );
  OR2 r253_U196 ( .A(r253_n40), .B(U3_U14_Z_7), .Z(r253_n41) );
  AO2 r253_U195 ( .A(U3_U14_Z_7), .B(r253_n40), .C(r253_n41), .D(U3_U18_Z_29), 
        .Z(r253_n38) );
  EO r253_U194 ( .A(r253_n37), .B(U3_U18_Z_30), .Z(r253_n39) );
  EO r253_U193 ( .A(r253_n38), .B(r253_n39), .Z(n287) );
  EO r253_U192 ( .A(U3_U18_Z_31), .B(r253_n37), .Z(r253_n34) );
  NR2 r253_U191 ( .A(r253_n38), .B(r253_n37), .Z(r253_n36) );
  EON1 r253_U190 ( .A(U3_U18_Z_30), .B(r253_n36), .C(r253_n37), .D(r253_n38), 
        .Z(r253_n35) );
  EO r253_U189 ( .A(r253_n34), .B(r253_n35), .Z(n286) );
  EO r253_U188 ( .A(U3_U18_Z_3), .B(r253_n33), .Z(r253_n32) );
  EO r253_U187 ( .A(r253_n25), .B(r253_n32), .Z(n314) );
  AN2 r253_U186 ( .A(r253_n29), .B(r253_n28), .Z(r253_n30) );
  AO4 r253_U185 ( .A(r253_n28), .B(r253_n29), .C(r253_n30), .D(r253_n31), .Z(
        r253_n26) );
  AN2 r253_U184 ( .A(r253_n26), .B(r253_n25), .Z(r253_n27) );
  AO4 r253_U183 ( .A(r253_n25), .B(r253_n26), .C(U3_U18_Z_3), .D(r253_n27), 
        .Z(r253_n17) );
  IV r253_U182 ( .A(U3_U18_Z_4), .Z(r253_n19) );
  EO r253_U181 ( .A(r253_n17), .B(r253_n19), .Z(r253_n24) );
  EN r253_U180 ( .A(r253_n16), .B(r253_n24), .Z(n313) );
  IV r253_U179 ( .A(r253_n23), .Z(r253_n13) );
  EO r253_U178 ( .A(r253_n21), .B(r253_n22), .Z(r253_n20) );
  EO r253_U177 ( .A(r253_n13), .B(r253_n20), .Z(n312) );
  AN2 r253_U176 ( .A(r253_n17), .B(r253_n16), .Z(r253_n18) );
  AO4 r253_U175 ( .A(r253_n16), .B(r253_n17), .C(r253_n18), .D(r253_n19), .Z(
        r253_n14) );
  AN2 r253_U174 ( .A(r253_n14), .B(r253_n13), .Z(r253_n15) );
  AO4 r253_U173 ( .A(r253_n13), .B(r253_n14), .C(U3_U18_Z_5), .D(r253_n15), 
        .Z(r253_n12) );
  EN r253_U172 ( .A(r253_n12), .B(U3_U18_Z_6), .Z(r253_n11) );
  EO r253_U171 ( .A(r253_n10), .B(r253_n11), .Z(n311) );
  EN r253_U170 ( .A(r253_n9), .B(U3_U18_Z_7), .Z(r253_n8) );
  EN r253_U169 ( .A(r253_n7), .B(r253_n8), .Z(n310) );
  EO r253_U168 ( .A(U3_U14_Z_7), .B(r253_n6), .Z(r253_n5) );
  EO r253_U167 ( .A(r253_n4), .B(r253_n5), .Z(n309) );
  EO r253_U166 ( .A(U3_U14_Z_7), .B(r253_n3), .Z(r253_n1) );
  EO r253_U165 ( .A(r253_n1), .B(r253_n2), .Z(n308) );
  EO r1161_U60 ( .A(U3_U4_Z_0), .B(U3_U3_Z_0), .Z(N1750) );
  AN3 r1161_U59 ( .A(U3_U3_Z_1), .B(U3_U3_Z_0), .C(U3_U4_Z_0), .Z(r1161_n8) );
  AN3 r1161_U58 ( .A(U3_U3_Z_2), .B(r1161_n8), .C(U3_U3_Z_3), .Z(r1161_n6) );
  AN3 r1161_U57 ( .A(U3_U3_Z_4), .B(r1161_n6), .C(U3_U3_Z_5), .Z(r1161_n4) );
  AN3 r1161_U56 ( .A(U3_U3_Z_6), .B(r1161_n4), .C(U3_U3_Z_7), .Z(r1161_n2) );
  AN3 r1161_U55 ( .A(U3_U3_Z_8), .B(r1161_n2), .C(U3_U3_Z_9), .Z(r1161_n14) );
  EO r1161_U54 ( .A(r1161_n14), .B(U3_U3_Z_10), .Z(N1760) );
  ND2 r1161_U53 ( .A(U3_U3_Z_10), .B(r1161_n14), .Z(r1161_n15) );
  EN r1161_U52 ( .A(r1161_n15), .B(U3_U3_Z_11), .Z(N1761) );
  AN3 r1161_U51 ( .A(U3_U3_Z_10), .B(r1161_n14), .C(U3_U3_Z_11), .Z(r1161_n13)
         );
  EO r1161_U50 ( .A(r1161_n13), .B(U3_U3_Z_12), .Z(N1762) );
  ND2 r1161_U49 ( .A(U3_U3_Z_12), .B(r1161_n13), .Z(r1161_n11) );
  EN r1161_U48 ( .A(r1161_n11), .B(U3_U3_Z_13), .Z(N1763) );
  IV r1161_U47 ( .A(U3_U3_Z_13), .Z(r1161_n12) );
  NR2 r1161_U46 ( .A(r1161_n11), .B(r1161_n12), .Z(r1161_n10) );
  EO r1161_U45 ( .A(U3_U3_Z_14), .B(r1161_n10), .Z(N1764) );
  ND2 r1161_U44 ( .A(U3_U4_Z_0), .B(U3_U3_Z_0), .Z(r1161_n9) );
  EN r1161_U43 ( .A(r1161_n9), .B(U3_U3_Z_1), .Z(N1751) );
  EO r1161_U42 ( .A(r1161_n8), .B(U3_U3_Z_2), .Z(N1752) );
  ND2 r1161_U41 ( .A(U3_U3_Z_2), .B(r1161_n8), .Z(r1161_n7) );
  EN r1161_U40 ( .A(r1161_n7), .B(U3_U3_Z_3), .Z(N1753) );
  EO r1161_U39 ( .A(r1161_n6), .B(U3_U3_Z_4), .Z(N1754) );
  ND2 r1161_U38 ( .A(U3_U3_Z_4), .B(r1161_n6), .Z(r1161_n5) );
  EN r1161_U37 ( .A(r1161_n5), .B(U3_U3_Z_5), .Z(N1755) );
  EO r1161_U36 ( .A(r1161_n4), .B(U3_U3_Z_6), .Z(N1756) );
  ND2 r1161_U35 ( .A(U3_U3_Z_6), .B(r1161_n4), .Z(r1161_n3) );
  EN r1161_U34 ( .A(r1161_n3), .B(U3_U3_Z_7), .Z(N1757) );
  EO r1161_U33 ( .A(r1161_n2), .B(U3_U3_Z_8), .Z(N1758) );
  ND2 r1161_U32 ( .A(U3_U3_Z_8), .B(r1161_n2), .Z(r1161_n1) );
  EN r1161_U31 ( .A(r1161_n1), .B(U3_U3_Z_9), .Z(N1759) );
  EO r1158_U183 ( .A(U3_U14_Z_7), .B(U3_U14_Z_0), .Z(r1158_n56) );
  EO r1158_U182 ( .A(U3_U13_Z_0), .B(r1158_n56), .Z(n460) );
  AO5 r1158_U181 ( .A(U3_U14_Z_0), .B(U3_U14_Z_7), .C(U3_U13_Z_0), .Z(
        r1158_n55) );
  IV r1158_U180 ( .A(r1158_n55), .Z(r1158_n30) );
  OR2 r1158_U179 ( .A(r1158_n30), .B(U3_U13_Z_1), .Z(r1158_n54) );
  AO2 r1158_U178 ( .A(r1158_n30), .B(U3_U13_Z_1), .C(r1158_n54), .D(U3_U14_Z_1), .Z(r1158_n18) );
  IV r1158_U177 ( .A(r1158_n18), .Z(r1158_n52) );
  OR2 r1158_U176 ( .A(U3_U13_Z_2), .B(r1158_n52), .Z(r1158_n53) );
  AO2 r1158_U175 ( .A(r1158_n52), .B(U3_U13_Z_2), .C(r1158_n53), .D(U3_U14_Z_2), .Z(r1158_n12) );
  IV r1158_U174 ( .A(r1158_n12), .Z(r1158_n50) );
  AN2 r1158_U173 ( .A(r1158_n50), .B(U3_U13_Z_3), .Z(r1158_n51) );
  AO4 r1158_U172 ( .A(U3_U13_Z_3), .B(r1158_n50), .C(U3_U14_Z_3), .D(r1158_n51), .Z(r1158_n11) );
  IV r1158_U171 ( .A(r1158_n11), .Z(r1158_n48) );
  OR2 r1158_U170 ( .A(r1158_n48), .B(U3_U13_Z_4), .Z(r1158_n49) );
  AO2 r1158_U169 ( .A(r1158_n48), .B(U3_U13_Z_4), .C(r1158_n49), .D(U3_U14_Z_4), .Z(r1158_n8) );
  IV r1158_U168 ( .A(r1158_n8), .Z(r1158_n46) );
  AN2 r1158_U167 ( .A(r1158_n46), .B(U3_U13_Z_5), .Z(r1158_n47) );
  AO4 r1158_U166 ( .A(U3_U13_Z_5), .B(r1158_n46), .C(U3_U14_Z_5), .D(r1158_n47), .Z(r1158_n7) );
  IV r1158_U165 ( .A(r1158_n7), .Z(r1158_n44) );
  OR2 r1158_U164 ( .A(r1158_n44), .B(U3_U13_Z_6), .Z(r1158_n45) );
  AO2 r1158_U163 ( .A(r1158_n44), .B(U3_U13_Z_6), .C(r1158_n45), .D(U3_U14_Z_6), .Z(r1158_n4) );
  IV r1158_U162 ( .A(r1158_n4), .Z(r1158_n42) );
  AN2 r1158_U161 ( .A(r1158_n42), .B(U3_U13_Z_7), .Z(r1158_n43) );
  AO4 r1158_U160 ( .A(U3_U13_Z_7), .B(r1158_n42), .C(U3_U14_Z_7), .D(r1158_n43), .Z(r1158_n2) );
  IV r1158_U159 ( .A(r1158_n2), .Z(r1158_n41) );
  AN3 r1158_U158 ( .A(r1158_n41), .B(U3_U13_Z_8), .C(U3_U13_Z_9), .Z(r1158_n39) );
  EO r1158_U157 ( .A(r1158_n39), .B(U3_U13_Z_10), .Z(n450) );
  ND2 r1158_U156 ( .A(U3_U13_Z_10), .B(r1158_n39), .Z(r1158_n40) );
  EN r1158_U155 ( .A(r1158_n40), .B(U3_U13_Z_11), .Z(n449) );
  AN3 r1158_U154 ( .A(U3_U13_Z_10), .B(r1158_n39), .C(U3_U13_Z_11), .Z(
        r1158_n37) );
  EO r1158_U153 ( .A(r1158_n37), .B(U3_U13_Z_12), .Z(n448) );
  ND2 r1158_U152 ( .A(U3_U13_Z_12), .B(r1158_n37), .Z(r1158_n38) );
  EN r1158_U151 ( .A(r1158_n38), .B(U3_U13_Z_13), .Z(n447) );
  AN3 r1158_U150 ( .A(U3_U13_Z_12), .B(r1158_n37), .C(U3_U13_Z_13), .Z(
        r1158_n35) );
  EO r1158_U149 ( .A(r1158_n35), .B(U3_U13_Z_14), .Z(n446) );
  ND2 r1158_U148 ( .A(U3_U13_Z_14), .B(r1158_n35), .Z(r1158_n36) );
  EN r1158_U147 ( .A(r1158_n36), .B(U3_U13_Z_15), .Z(n445) );
  AN3 r1158_U146 ( .A(U3_U13_Z_14), .B(r1158_n35), .C(U3_U13_Z_15), .Z(
        r1158_n33) );
  EO r1158_U145 ( .A(r1158_n33), .B(U3_U13_Z_16), .Z(n444) );
  ND2 r1158_U144 ( .A(U3_U13_Z_16), .B(r1158_n33), .Z(r1158_n34) );
  EN r1158_U143 ( .A(r1158_n34), .B(U3_U13_Z_17), .Z(n443) );
  AN3 r1158_U142 ( .A(U3_U13_Z_16), .B(r1158_n33), .C(U3_U13_Z_17), .Z(
        r1158_n29) );
  EO r1158_U141 ( .A(r1158_n29), .B(U3_U13_Z_18), .Z(n442) );
  ND2 r1158_U140 ( .A(U3_U13_Z_18), .B(r1158_n29), .Z(r1158_n32) );
  EN r1158_U139 ( .A(r1158_n32), .B(U3_U13_Z_19), .Z(n441) );
  EO r1158_U138 ( .A(U3_U14_Z_1), .B(U3_U13_Z_1), .Z(r1158_n31) );
  EO r1158_U137 ( .A(r1158_n30), .B(r1158_n31), .Z(n459) );
  AN3 r1158_U136 ( .A(U3_U13_Z_18), .B(r1158_n29), .C(U3_U13_Z_19), .Z(
        r1158_n27) );
  EO r1158_U135 ( .A(r1158_n27), .B(U3_U13_Z_20), .Z(n440) );
  ND2 r1158_U134 ( .A(U3_U13_Z_20), .B(r1158_n27), .Z(r1158_n28) );
  EN r1158_U133 ( .A(r1158_n28), .B(U3_U13_Z_21), .Z(n439) );
  AN3 r1158_U132 ( .A(U3_U13_Z_20), .B(r1158_n27), .C(U3_U13_Z_21), .Z(
        r1158_n25) );
  EO r1158_U131 ( .A(r1158_n25), .B(U3_U13_Z_22), .Z(n438) );
  ND2 r1158_U130 ( .A(U3_U13_Z_22), .B(r1158_n25), .Z(r1158_n26) );
  EN r1158_U129 ( .A(r1158_n26), .B(U3_U13_Z_23), .Z(n437) );
  AN3 r1158_U128 ( .A(U3_U13_Z_22), .B(r1158_n25), .C(U3_U13_Z_23), .Z(
        r1158_n23) );
  EO r1158_U127 ( .A(r1158_n23), .B(U3_U13_Z_24), .Z(n436) );
  ND2 r1158_U126 ( .A(U3_U13_Z_24), .B(r1158_n23), .Z(r1158_n24) );
  EN r1158_U125 ( .A(r1158_n24), .B(U3_U13_Z_25), .Z(n435) );
  AN3 r1158_U124 ( .A(U3_U13_Z_24), .B(r1158_n23), .C(U3_U13_Z_25), .Z(
        r1158_n21) );
  EO r1158_U123 ( .A(r1158_n21), .B(U3_U13_Z_26), .Z(n434) );
  ND2 r1158_U122 ( .A(U3_U13_Z_26), .B(r1158_n21), .Z(r1158_n22) );
  EN r1158_U121 ( .A(r1158_n22), .B(U3_U13_Z_27), .Z(n433) );
  AN3 r1158_U120 ( .A(U3_U13_Z_26), .B(r1158_n21), .C(U3_U13_Z_27), .Z(
        r1158_n20) );
  EO r1158_U119 ( .A(r1158_n20), .B(U3_U13_Z_28), .Z(n432) );
  AN2 r1158_U118 ( .A(U3_U13_Z_28), .B(r1158_n20), .Z(r1158_n17) );
  EO r1158_U117 ( .A(r1158_n17), .B(U3_U13_Z_29), .Z(n431) );
  EN r1158_U116 ( .A(U3_U14_Z_2), .B(U3_U13_Z_2), .Z(r1158_n19) );
  EO r1158_U115 ( .A(r1158_n18), .B(r1158_n19), .Z(n458) );
  ND2 r1158_U114 ( .A(U3_U13_Z_29), .B(r1158_n17), .Z(r1158_n15) );
  IV r1158_U113 ( .A(U3_U13_Z_30), .Z(r1158_n16) );
  EO r1158_U112 ( .A(r1158_n15), .B(r1158_n16), .Z(n430) );
  NR2 r1158_U111 ( .A(r1158_n15), .B(r1158_n16), .Z(r1158_n14) );
  EO r1158_U110 ( .A(U3_U13_Z_31), .B(r1158_n14), .Z(n429) );
  EN r1158_U109 ( .A(U3_U14_Z_3), .B(U3_U13_Z_3), .Z(r1158_n13) );
  EO r1158_U108 ( .A(r1158_n12), .B(r1158_n13), .Z(n457) );
  EN r1158_U107 ( .A(U3_U14_Z_4), .B(U3_U13_Z_4), .Z(r1158_n10) );
  EO r1158_U106 ( .A(r1158_n10), .B(r1158_n11), .Z(n456) );
  EN r1158_U105 ( .A(U3_U14_Z_5), .B(U3_U13_Z_5), .Z(r1158_n9) );
  EO r1158_U104 ( .A(r1158_n8), .B(r1158_n9), .Z(n455) );
  EN r1158_U103 ( .A(U3_U14_Z_6), .B(U3_U13_Z_6), .Z(r1158_n6) );
  EO r1158_U102 ( .A(r1158_n6), .B(r1158_n7), .Z(n454) );
  EN r1158_U101 ( .A(U3_U14_Z_7), .B(U3_U13_Z_7), .Z(r1158_n5) );
  EO r1158_U100 ( .A(r1158_n4), .B(r1158_n5), .Z(n453) );
  IV r1158_U99 ( .A(U3_U13_Z_8), .Z(r1158_n3) );
  EO r1158_U98 ( .A(r1158_n2), .B(r1158_n3), .Z(n452) );
  NR2 r1158_U97 ( .A(r1158_n2), .B(r1158_n3), .Z(r1158_n1) );
  EO r1158_U96 ( .A(U3_U13_Z_9), .B(r1158_n1), .Z(n451) );
  EO r1160_U121 ( .A(U3_U1_Z_0), .B(U3_U2_Z_0), .Z(N558) );
  AN3 r1160_U120 ( .A(U3_U1_Z_0), .B(U3_U2_Z_0), .C(U3_U1_Z_1), .Z(r1160_n9)
         );
  AN3 r1160_U119 ( .A(U3_U1_Z_2), .B(r1160_n9), .C(U3_U1_Z_3), .Z(r1160_n7) );
  AN3 r1160_U118 ( .A(U3_U1_Z_4), .B(r1160_n7), .C(U3_U1_Z_5), .Z(r1160_n5) );
  AN3 r1160_U117 ( .A(U3_U1_Z_6), .B(r1160_n5), .C(U3_U1_Z_7), .Z(r1160_n3) );
  AN3 r1160_U116 ( .A(U3_U1_Z_8), .B(r1160_n3), .C(U3_U1_Z_9), .Z(r1160_n29)
         );
  EO r1160_U115 ( .A(r1160_n29), .B(U3_U1_Z_10), .Z(N568) );
  ND2 r1160_U114 ( .A(U3_U1_Z_10), .B(r1160_n29), .Z(r1160_n30) );
  EN r1160_U113 ( .A(r1160_n30), .B(U3_U1_Z_11), .Z(N569) );
  AN3 r1160_U112 ( .A(U3_U1_Z_10), .B(r1160_n29), .C(U3_U1_Z_11), .Z(r1160_n27) );
  EO r1160_U111 ( .A(r1160_n27), .B(U3_U1_Z_12), .Z(N570) );
  ND2 r1160_U110 ( .A(U3_U1_Z_12), .B(r1160_n27), .Z(r1160_n28) );
  EN r1160_U109 ( .A(r1160_n28), .B(U3_U1_Z_13), .Z(N571) );
  AN3 r1160_U108 ( .A(U3_U1_Z_12), .B(r1160_n27), .C(U3_U1_Z_13), .Z(r1160_n25) );
  EO r1160_U107 ( .A(r1160_n25), .B(U3_U1_Z_14), .Z(N572) );
  ND2 r1160_U106 ( .A(U3_U1_Z_14), .B(r1160_n25), .Z(r1160_n26) );
  EN r1160_U105 ( .A(r1160_n26), .B(U3_U1_Z_15), .Z(N573) );
  AN3 r1160_U104 ( .A(U3_U1_Z_14), .B(r1160_n25), .C(U3_U1_Z_15), .Z(r1160_n23) );
  EO r1160_U103 ( .A(r1160_n23), .B(U3_U1_Z_16), .Z(N574) );
  ND2 r1160_U102 ( .A(U3_U1_Z_16), .B(r1160_n23), .Z(r1160_n24) );
  EN r1160_U101 ( .A(r1160_n24), .B(U3_U1_Z_17), .Z(N575) );
  AN3 r1160_U100 ( .A(U3_U1_Z_16), .B(r1160_n23), .C(U3_U1_Z_17), .Z(r1160_n20) );
  EO r1160_U99 ( .A(r1160_n20), .B(U3_U1_Z_18), .Z(N576) );
  ND2 r1160_U98 ( .A(U3_U1_Z_18), .B(r1160_n20), .Z(r1160_n22) );
  EN r1160_U97 ( .A(r1160_n22), .B(U3_U1_Z_19), .Z(N577) );
  ND2 r1160_U96 ( .A(U3_U1_Z_0), .B(U3_U2_Z_0), .Z(r1160_n21) );
  EN r1160_U95 ( .A(r1160_n21), .B(U3_U1_Z_1), .Z(N559) );
  AN3 r1160_U94 ( .A(U3_U1_Z_18), .B(r1160_n20), .C(U3_U1_Z_19), .Z(r1160_n18)
         );
  EO r1160_U93 ( .A(r1160_n18), .B(U3_U1_Z_20), .Z(N578) );
  ND2 r1160_U92 ( .A(U3_U1_Z_20), .B(r1160_n18), .Z(r1160_n19) );
  EN r1160_U91 ( .A(r1160_n19), .B(U3_U1_Z_21), .Z(N579) );
  AN3 r1160_U90 ( .A(U3_U1_Z_20), .B(r1160_n18), .C(U3_U1_Z_21), .Z(r1160_n16)
         );
  EO r1160_U89 ( .A(r1160_n16), .B(U3_U1_Z_22), .Z(N580) );
  ND2 r1160_U88 ( .A(U3_U1_Z_22), .B(r1160_n16), .Z(r1160_n17) );
  EN r1160_U87 ( .A(r1160_n17), .B(U3_U1_Z_23), .Z(N581) );
  AN3 r1160_U86 ( .A(U3_U1_Z_22), .B(r1160_n16), .C(U3_U1_Z_23), .Z(r1160_n14)
         );
  EO r1160_U85 ( .A(r1160_n14), .B(U3_U1_Z_24), .Z(N582) );
  ND2 r1160_U84 ( .A(U3_U1_Z_24), .B(r1160_n14), .Z(r1160_n15) );
  EN r1160_U83 ( .A(r1160_n15), .B(U3_U1_Z_25), .Z(N583) );
  AN3 r1160_U82 ( .A(U3_U1_Z_24), .B(r1160_n14), .C(U3_U1_Z_25), .Z(r1160_n13)
         );
  EO r1160_U81 ( .A(r1160_n13), .B(U3_U1_Z_26), .Z(N584) );
  EO r1160_U80 ( .A(r1160_n1), .B(U3_U1_Z_27), .Z(N585) );
  ND2 r1160_U79 ( .A(U3_U1_Z_27), .B(r1160_n1), .Z(r1160_n11) );
  EN r1160_U78 ( .A(r1160_n11), .B(U3_U1_Z_28), .Z(N586) );
  IV r1160_U77 ( .A(U3_U1_Z_28), .Z(r1160_n12) );
  NR2 r1160_U76 ( .A(r1160_n11), .B(r1160_n12), .Z(r1160_n10) );
  EO r1160_U75 ( .A(U3_U1_Z_29), .B(r1160_n10), .Z(N587) );
  EO r1160_U74 ( .A(r1160_n9), .B(U3_U1_Z_2), .Z(N560) );
  ND2 r1160_U73 ( .A(U3_U1_Z_2), .B(r1160_n9), .Z(r1160_n8) );
  EN r1160_U72 ( .A(r1160_n8), .B(U3_U1_Z_3), .Z(N561) );
  EO r1160_U71 ( .A(r1160_n7), .B(U3_U1_Z_4), .Z(N562) );
  ND2 r1160_U70 ( .A(U3_U1_Z_4), .B(r1160_n7), .Z(r1160_n6) );
  EN r1160_U69 ( .A(r1160_n6), .B(U3_U1_Z_5), .Z(N563) );
  EO r1160_U68 ( .A(r1160_n5), .B(U3_U1_Z_6), .Z(N564) );
  ND2 r1160_U67 ( .A(U3_U1_Z_6), .B(r1160_n5), .Z(r1160_n4) );
  EN r1160_U66 ( .A(r1160_n4), .B(U3_U1_Z_7), .Z(N565) );
  EO r1160_U65 ( .A(r1160_n3), .B(U3_U1_Z_8), .Z(N566) );
  ND2 r1160_U64 ( .A(U3_U1_Z_8), .B(r1160_n3), .Z(r1160_n2) );
  EN r1160_U63 ( .A(r1160_n2), .B(U3_U1_Z_9), .Z(N567) );
  AN2I r1160_U62 ( .A(U3_U1_Z_26), .B(r1160_n13), .Z(r1160_n1) );
endmodule

